task test_rectangle();
    $display("RECTANGLE Program");
endtask