task test_ctr_aes();
    $display("CTR AES Program");
endtask