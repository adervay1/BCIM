// avalon_mm_sim_block.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module avalon_mm_sim_block (
		input  wire        clk,               //       clk.clk
		input  wire        reset,             // clk_reset.reset
		output wire [31:0] avm_address,       //        m0.address
		input  wire [31:0] avm_readdata,      //          .readdata
		output wire [31:0] avm_writedata,     //          .writedata
		input  wire        avm_waitrequest,   //          .waitrequest
		output wire        avm_write,         //          .write
		output wire        avm_read,          //          .read
		input  wire        avm_readdatavalid  //          .readdatavalid
	);

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (32),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (4),
		.AV_BURSTCOUNT_W            (1),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (0),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (1),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (0)
	) mm_master_bfm_0 (
		.clk                    (clk),               //       clk.clk
		.reset                  (reset),             // clk_reset.reset
		.avm_address            (avm_address),       //        m0.address
		.avm_readdata           (avm_readdata),      //          .readdata
		.avm_writedata          (avm_writedata),     //          .writedata
		.avm_waitrequest        (avm_waitrequest),   //          .waitrequest
		.avm_write              (avm_write),         //          .write
		.avm_read               (avm_read),          //          .read
		.avm_readdatavalid      (avm_readdatavalid), //          .readdatavalid
		.avm_burstcount         (),                  // (terminated)
		.avm_begintransfer      (),                  // (terminated)
		.avm_beginbursttransfer (),                  // (terminated)
		.avm_byteenable         (),                  // (terminated)
		.avm_arbiterlock        (),                  // (terminated)
		.avm_lock               (),                  // (terminated)
		.avm_debugaccess        (),                  // (terminated)
		.avm_transactionid      (),                  // (terminated)
		.avm_readid             (8'b00000000),       // (terminated)
		.avm_writeid            (8'b00000000),       // (terminated)
		.avm_clken              (),                  // (terminated)
		.avm_response           (2'b00),             // (terminated)
		.avm_writeresponsevalid (1'b0),              // (terminated)
		.avm_readresponse       (8'b00000000),       // (terminated)
		.avm_writeresponse      (8'b00000000)        // (terminated)
	);

endmodule
