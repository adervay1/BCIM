//TODO: Delete
task test_ecb_aes();
    $display("ECB AES Program");
endtask

//Rounds
task AES_ECB_Encrypt();
    logic [7:0] state_bytes [15:0];
    logic [7:0] plain_text_bytes [15:0];
    logic [7:0] round_key_bytes [15:0];
    logic [7:0] key_bytes [9:0][15:0];

    //Load Plain Text
    //Column-Wise 0-3
    plain_text_bytes    = '{8'h32,8'h88,8'h31,8'hE0,  //Row 0
                            8'h43,8'h5A,8'h31,8'h37,
                            8'hF6,8'h30,8'h98,8'h07,
                            8'hA8,8'h8D,8'hA2,8'h34}; //Row 3
    Load_AES_State_1Col(plain_text_bytes,'h0);
    
    //#10us;
    //Print_State_Bytes_1Col('h0,"Plain Text:");
    
    
    round_key_bytes = '{8'h2B,8'h28,8'hAB,8'h09,  //Row 0
                        8'h7E,8'hAE,8'hF7,8'hCF,
                        8'h15,8'hD2,8'h15,8'h4F,
                        8'h16,8'hA6,8'h88,8'h3C}; //Row 3
    Load_AES_State_1Col(round_key_bytes,'h80);
    
    //#10us;
    //Print_State_Bytes_1Col('h80,"Initial Key");
    
    AES_ARK();
    
    //#10us;
    //Print_State_Bytes_1Col('h00,"Initial Add Key");
    
    
    
    AES_SBOX();
    
    //#10us;
    //Print_State_Bytes_1Col('h00,"Initial Add Key");
    
    AES_MC();
    
    //#10us;
    //Print_State_Bytes_1Col('h80,"1 Col");
    
    
    
    key_bytes[0] = '{8'hA0,8'h88,8'h23,8'h2A,  //Row 0
                    8'hFA,8'h54,8'hA3,8'h6C,
                    8'hFE,8'h2C,8'h39,8'h76,
                    8'h17,8'hB1,8'h39,8'h05}; //Row 3
    Load_AES_State_1Col(key_bytes[0],'h00);
    
    
    AES_ARK();
    
    #10us;
    Print_AES_State_Bytes_1Col('h00,"Add Key 1");

endtask


task AES_ECB_Decrypt();
    logic [7:0] round_key_bytes [15:0];
    logic [7:0] key_bytes [9:0][15:0];

    key_bytes[0] = '{8'hA0,8'h88,8'h23,8'h2A,  //Row 0
                    8'hFA,8'h54,8'hA3,8'h6C,
                    8'hFE,8'h2C,8'h39,8'h76,
                    8'h17,8'hB1,8'h39,8'h05}; //Row 3
    Load_AES_State_1Col(key_bytes[0],'h80);
    
    
    AES_ARK();
    
    #10us;
    Print_AES_State_Bytes_1Col('h00,"Inv Add Key 1");
    
    
    AES_Inv_MC();
    
    #10us;
    Print_AES_State_Bytes_1Col('h80,"Inv Mix Cols");
    
    
    AES_Inv_SBOX();
    
    #10us;
    Print_AES_State_Bytes_1Col('h80,"Inv SBOX");
    
    round_key_bytes = '{8'h2B,8'h28,8'hAB,8'h09,  //Row 0
                        8'h7E,8'hAE,8'hF7,8'hCF,
                        8'h15,8'hD2,8'h15,8'h4F,
                        8'h16,8'hA6,8'h88,8'h3C}; //Row 3
    Load_AES_State_1Col(round_key_bytes,'h00);
    
    
    AES_ARK();
    
    #10us;
    Print_AES_State_Bytes_1Col('h00,"Plaintext");


endtask


//Common / Utility
task Load_AES_State_1Col(input logic [7:0] byte_in [15:0], input int start_addr);
    Load_IMC_Byte(byte_in[15],start_addr+'h0);
    Load_IMC_Byte(byte_in[11],start_addr+'h8);
    Load_IMC_Byte(byte_in[7],start_addr+'h10);
    Load_IMC_Byte(byte_in[3],start_addr+'h18);

    Load_IMC_Byte(byte_in[14],start_addr+'h20);
    Load_IMC_Byte(byte_in[10],start_addr+'h28);
    Load_IMC_Byte(byte_in[6],start_addr+'h30);
    Load_IMC_Byte(byte_in[2],start_addr+'h38);

    Load_IMC_Byte(byte_in[13],start_addr+'h40);
    Load_IMC_Byte(byte_in[9],start_addr+'h48);
    Load_IMC_Byte(byte_in[5],start_addr+'h50);
    Load_IMC_Byte(byte_in[1],start_addr+'h58);

    Load_IMC_Byte(byte_in[12],start_addr+'h60);
    Load_IMC_Byte(byte_in[8],start_addr+'h68);
    Load_IMC_Byte(byte_in[4],start_addr+'h70);
    Load_IMC_Byte(byte_in[0],start_addr+'h78);
endtask


//Round Functions

task AES_ARK();
//State Input   00-7F
//Key Input     80-FF
//Output        00-7F

    Send_IMC_Command(32'd83918848);
    Send_IMC_Command(32'd83984641);
    Send_IMC_Command(32'd84050434);
    Send_IMC_Command(32'd84116227);
    Send_IMC_Command(32'd84182020);
    Send_IMC_Command(32'd84247813);
    Send_IMC_Command(32'd84313606);
    Send_IMC_Command(32'd84379399);
    Send_IMC_Command(32'd84445192);
    Send_IMC_Command(32'd84510985);
    Send_IMC_Command(32'd84576778);
    Send_IMC_Command(32'd84642571);
    Send_IMC_Command(32'd84708364);
    Send_IMC_Command(32'd84774157);
    Send_IMC_Command(32'd84839950);
    Send_IMC_Command(32'd84905743);
    Send_IMC_Command(32'd84971536);
    Send_IMC_Command(32'd85037329);
    Send_IMC_Command(32'd85103122);
    Send_IMC_Command(32'd85168915);
    Send_IMC_Command(32'd85234708);
    Send_IMC_Command(32'd85300501);
    Send_IMC_Command(32'd85366294);
    Send_IMC_Command(32'd85432087);
    Send_IMC_Command(32'd85497880);
    Send_IMC_Command(32'd85563673);
    Send_IMC_Command(32'd85629466);
    Send_IMC_Command(32'd85695259);
    Send_IMC_Command(32'd85761052);
    Send_IMC_Command(32'd85826845);
    Send_IMC_Command(32'd85892638);
    Send_IMC_Command(32'd85958431);
    Send_IMC_Command(32'd86024224);
    Send_IMC_Command(32'd86090017);
    Send_IMC_Command(32'd86155810);
    Send_IMC_Command(32'd86221603);
    Send_IMC_Command(32'd86287396);
    Send_IMC_Command(32'd86353189);
    Send_IMC_Command(32'd86418982);
    Send_IMC_Command(32'd86484775);
    Send_IMC_Command(32'd86550568);
    Send_IMC_Command(32'd86616361);
    Send_IMC_Command(32'd86682154);
    Send_IMC_Command(32'd86747947);
    Send_IMC_Command(32'd86813740);
    Send_IMC_Command(32'd86879533);
    Send_IMC_Command(32'd86945326);
    Send_IMC_Command(32'd87011119);
    Send_IMC_Command(32'd87076912);
    Send_IMC_Command(32'd87142705);
    Send_IMC_Command(32'd87208498);
    Send_IMC_Command(32'd87274291);
    Send_IMC_Command(32'd87340084);
    Send_IMC_Command(32'd87405877);
    Send_IMC_Command(32'd87471670);
    Send_IMC_Command(32'd87537463);
    Send_IMC_Command(32'd87603256);
    Send_IMC_Command(32'd87669049);
    Send_IMC_Command(32'd87734842);
    Send_IMC_Command(32'd87800635);
    Send_IMC_Command(32'd87866428);
    Send_IMC_Command(32'd87932221);
    Send_IMC_Command(32'd87998014);
    Send_IMC_Command(32'd88063807);
    Send_IMC_Command(32'd88129600);
    Send_IMC_Command(32'd88195393);
    Send_IMC_Command(32'd88261186);
    Send_IMC_Command(32'd88326979);
    Send_IMC_Command(32'd88392772);
    Send_IMC_Command(32'd88458565);
    Send_IMC_Command(32'd88524358);
    Send_IMC_Command(32'd88590151);
    Send_IMC_Command(32'd88655944);
    Send_IMC_Command(32'd88721737);
    Send_IMC_Command(32'd88787530);
    Send_IMC_Command(32'd88853323);
    Send_IMC_Command(32'd88919116);
    Send_IMC_Command(32'd88984909);
    Send_IMC_Command(32'd89050702);
    Send_IMC_Command(32'd89116495);
    Send_IMC_Command(32'd89182288);
    Send_IMC_Command(32'd89248081);
    Send_IMC_Command(32'd89313874);
    Send_IMC_Command(32'd89379667);
    Send_IMC_Command(32'd89445460);
    Send_IMC_Command(32'd89511253);
    Send_IMC_Command(32'd89577046);
    Send_IMC_Command(32'd89642839);
    Send_IMC_Command(32'd89708632);
    Send_IMC_Command(32'd89774425);
    Send_IMC_Command(32'd89840218);
    Send_IMC_Command(32'd89906011);
    Send_IMC_Command(32'd89971804);
    Send_IMC_Command(32'd90037597);
    Send_IMC_Command(32'd90103390);
    Send_IMC_Command(32'd90169183);
    Send_IMC_Command(32'd90234976);
    Send_IMC_Command(32'd90300769);
    Send_IMC_Command(32'd90366562);
    Send_IMC_Command(32'd90432355);
    Send_IMC_Command(32'd90498148);
    Send_IMC_Command(32'd90563941);
    Send_IMC_Command(32'd90629734);
    Send_IMC_Command(32'd90695527);
    Send_IMC_Command(32'd90761320);
    Send_IMC_Command(32'd90827113);
    Send_IMC_Command(32'd90892906);
    Send_IMC_Command(32'd90958699);
    Send_IMC_Command(32'd91024492);
    Send_IMC_Command(32'd91090285);
    Send_IMC_Command(32'd91156078);
    Send_IMC_Command(32'd91221871);
    Send_IMC_Command(32'd91287664);
    Send_IMC_Command(32'd91353457);
    Send_IMC_Command(32'd91419250);
    Send_IMC_Command(32'd91485043);
    Send_IMC_Command(32'd91550836);
    Send_IMC_Command(32'd91616629);
    Send_IMC_Command(32'd91682422);
    Send_IMC_Command(32'd91748215);
    Send_IMC_Command(32'd91814008);
    Send_IMC_Command(32'd91879801);
    Send_IMC_Command(32'd91945594);
    Send_IMC_Command(32'd92011387);
    Send_IMC_Command(32'd92077180);
    Send_IMC_Command(32'd92142973);
    Send_IMC_Command(32'd92208766);
    Send_IMC_Command(32'd92274559);
endtask

task AES_SBOX();

    Send_IMC_Command(32'd84148864);
    Send_IMC_Command(32'd84345217);
    Send_IMC_Command(32'd84345986);
    Send_IMC_Command(32'd84345475);
    Send_IMC_Command(32'd84280725);
    Send_IMC_Command(32'd93651076);
    Send_IMC_Command(32'd92537989);
    Send_IMC_Command(32'd92373126);
    Send_IMC_Command(32'd92538759);
    Send_IMC_Command(32'd92537224);
    Send_IMC_Command(32'd92832649);
    Send_IMC_Command(32'd84117142);
    Send_IMC_Command(32'd93717130);
    Send_IMC_Command(32'd93718155);
    Send_IMC_Command(32'd92930188);
    Send_IMC_Command(32'd92968333);
    Send_IMC_Command(32'd93029006);
    Send_IMC_Command(32'd83922575);
    Send_IMC_Command(32'd93163152);
    Send_IMC_Command(32'd93160337);
    Send_IMC_Command(32'd93687442);
    Send_IMC_Command(32'd92377747);
    Send_IMC_Command(32'd84382356);
    Send_IMC_Command(32'd75926167);
    Send_IMC_Command(32'd76123288);
    Send_IMC_Command(32'd93886361);
    Send_IMC_Command(32'd75825306);
    Send_IMC_Command(32'd94017435);
    Send_IMC_Command(32'd75600540);
    Send_IMC_Command(32'd76055709);
    Send_IMC_Command(32'd94215326);
    Send_IMC_Command(32'd75992991);
    Send_IMC_Command(32'd94346400);
    Send_IMC_Command(32'd75665057);
    Send_IMC_Command(32'd75534498);
    Send_IMC_Command(32'd94544291);
    Send_IMC_Command(32'd75730340);
    Send_IMC_Command(32'd94675365);
    Send_IMC_Command(32'd93948838);
    Send_IMC_Command(32'd94086567);
    Send_IMC_Command(32'd94282664);
    Send_IMC_Command(32'd94414249);
    Send_IMC_Command(32'd94806954);
    Send_IMC_Command(32'd94867883);
    Send_IMC_Command(32'd94933932);
    Send_IMC_Command(32'd94999725);
    Send_IMC_Command(32'd95071150);
    Send_IMC_Command(32'd78294191);
    Send_IMC_Command(32'd95268784);
    Send_IMC_Command(32'd78557361);
    Send_IMC_Command(32'd95529906);
    Send_IMC_Command(32'd95202739);
    Send_IMC_Command(32'd95137716);
    Send_IMC_Command(32'd78951349);
    Send_IMC_Command(32'd95792566);
    Send_IMC_Command(32'd95205047);
    Send_IMC_Command(32'd95467192);
    Send_IMC_Command(32'd78493881);
    Send_IMC_Command(32'd96057274);
    Send_IMC_Command(32'd95467963);
    Send_IMC_Command(32'd78822332);
    Send_IMC_Command(32'd95337661);
    Send_IMC_Command(32'd96320190);
    Send_IMC_Command(32'd95598271);
    Send_IMC_Command(32'd95600064);
    Send_IMC_Command(32'd95861441);
    Send_IMC_Command(32'd96452290);
    Send_IMC_Command(32'd79792835);
    Send_IMC_Command(32'd79334596);
    Send_IMC_Command(32'd79036613);
    Send_IMC_Command(32'd79729350);
    Send_IMC_Command(32'd79529159);
    Send_IMC_Command(32'd78811080);
    Send_IMC_Command(32'd79662793);
    Send_IMC_Command(32'd79859914);
    Send_IMC_Command(32'd79597003);
    Send_IMC_Command(32'd79791820);
    Send_IMC_Command(32'd79333837);
    Send_IMC_Command(32'd79070670);
    Send_IMC_Command(32'd79725007);
    Send_IMC_Command(32'd79530192);
    Send_IMC_Command(32'd78809041);
    Send_IMC_Command(32'd79659730);
    Send_IMC_Command(32'd79855827);
    Send_IMC_Command(32'd79594452);
    Send_IMC_Command(32'd97702869);
    Send_IMC_Command(32'd97375702);
    Send_IMC_Command(32'd97310423);
    Send_IMC_Command(32'd96716248);
    Send_IMC_Command(32'd96781273);
    Send_IMC_Command(32'd96913370);
    Send_IMC_Command(32'd97507547);
    Send_IMC_Command(32'd97180380);
    Send_IMC_Command(32'd97246173);
    Send_IMC_Command(32'd98360798);
    Send_IMC_Command(32'd98228703);
    Send_IMC_Command(32'd96913632);
    Send_IMC_Command(32'd97572321);
    Send_IMC_Command(32'd98099426);
    Send_IMC_Command(32'd98033412);
    Send_IMC_Command(32'd97115363);
    Send_IMC_Command(32'd97640164);
    Send_IMC_Command(32'd98689765);
    Send_IMC_Command(32'd298837248);
    Send_IMC_Command(32'd97706982);
    Send_IMC_Command(32'd97963751);
    Send_IMC_Command(32'd98034439);
    Send_IMC_Command(32'd299820289);
    Send_IMC_Command(32'd98698243);
    Send_IMC_Command(32'd285532934);
    Send_IMC_Command(32'd98887400);
    Send_IMC_Command(32'd300471301);
    Send_IMC_Command(32'd99083266);
    Send_IMC_Command(32'd84675200);
    Send_IMC_Command(32'd84871553);
    Send_IMC_Command(32'd84872322);
    Send_IMC_Command(32'd84871811);
    Send_IMC_Command(32'd84807061);
    Send_IMC_Command(32'd93653124);
    Send_IMC_Command(32'd92540037);
    Send_IMC_Command(32'd92373126);
    Send_IMC_Command(32'd92540807);
    Send_IMC_Command(32'd92539272);
    Send_IMC_Command(32'd92832649);
    Send_IMC_Command(32'd84641430);
    Send_IMC_Command(32'd93719178);
    Send_IMC_Command(32'd93720203);
    Send_IMC_Command(32'd92932236);
    Send_IMC_Command(32'd92968333);
    Send_IMC_Command(32'd93029006);
    Send_IMC_Command(32'd84446863);
    Send_IMC_Command(32'd93163152);
    Send_IMC_Command(32'd93160337);
    Send_IMC_Command(32'd93687442);
    Send_IMC_Command(32'd92377747);
    Send_IMC_Command(32'd84906644);
    Send_IMC_Command(32'd75926167);
    Send_IMC_Command(32'd76123288);
    Send_IMC_Command(32'd93886361);
    Send_IMC_Command(32'd75827354);
    Send_IMC_Command(32'd94017435);
    Send_IMC_Command(32'd75600540);
    Send_IMC_Command(32'd76055709);
    Send_IMC_Command(32'd94215326);
    Send_IMC_Command(32'd75992991);
    Send_IMC_Command(32'd94346400);
    Send_IMC_Command(32'd75665057);
    Send_IMC_Command(32'd75534498);
    Send_IMC_Command(32'd94544291);
    Send_IMC_Command(32'd75730340);
    Send_IMC_Command(32'd94675365);
    Send_IMC_Command(32'd93948838);
    Send_IMC_Command(32'd94086567);
    Send_IMC_Command(32'd94282664);
    Send_IMC_Command(32'd94414249);
    Send_IMC_Command(32'd94806954);
    Send_IMC_Command(32'd94867883);
    Send_IMC_Command(32'd94933932);
    Send_IMC_Command(32'd94999725);
    Send_IMC_Command(32'd95071150);
    Send_IMC_Command(32'd78294191);
    Send_IMC_Command(32'd95268784);
    Send_IMC_Command(32'd78557361);
    Send_IMC_Command(32'd95529906);
    Send_IMC_Command(32'd95202739);
    Send_IMC_Command(32'd95137716);
    Send_IMC_Command(32'd78951349);
    Send_IMC_Command(32'd95792566);
    Send_IMC_Command(32'd95205047);
    Send_IMC_Command(32'd95467192);
    Send_IMC_Command(32'd78493881);
    Send_IMC_Command(32'd96057274);
    Send_IMC_Command(32'd95467963);
    Send_IMC_Command(32'd78822332);
    Send_IMC_Command(32'd95337661);
    Send_IMC_Command(32'd96320190);
    Send_IMC_Command(32'd95598271);
    Send_IMC_Command(32'd95600064);
    Send_IMC_Command(32'd95861441);
    Send_IMC_Command(32'd96452290);
    Send_IMC_Command(32'd79792835);
    Send_IMC_Command(32'd79334596);
    Send_IMC_Command(32'd79038661);
    Send_IMC_Command(32'd79729350);
    Send_IMC_Command(32'd79529159);
    Send_IMC_Command(32'd78811080);
    Send_IMC_Command(32'd79662793);
    Send_IMC_Command(32'd79859914);
    Send_IMC_Command(32'd79597003);
    Send_IMC_Command(32'd79791820);
    Send_IMC_Command(32'd79333837);
    Send_IMC_Command(32'd79070670);
    Send_IMC_Command(32'd79725007);
    Send_IMC_Command(32'd79530192);
    Send_IMC_Command(32'd78809041);
    Send_IMC_Command(32'd79659730);
    Send_IMC_Command(32'd79855827);
    Send_IMC_Command(32'd79594452);
    Send_IMC_Command(32'd97702869);
    Send_IMC_Command(32'd97375702);
    Send_IMC_Command(32'd97310423);
    Send_IMC_Command(32'd96716248);
    Send_IMC_Command(32'd96781273);
    Send_IMC_Command(32'd96913370);
    Send_IMC_Command(32'd97507547);
    Send_IMC_Command(32'd97180380);
    Send_IMC_Command(32'd97246173);
    Send_IMC_Command(32'd98360798);
    Send_IMC_Command(32'd98228703);
    Send_IMC_Command(32'd96913632);
    Send_IMC_Command(32'd97572321);
    Send_IMC_Command(32'd98099426);
    Send_IMC_Command(32'd98033420);
    Send_IMC_Command(32'd97115363);
    Send_IMC_Command(32'd97640164);
    Send_IMC_Command(32'd98689765);
    Send_IMC_Command(32'd298837256);
    Send_IMC_Command(32'd97706982);
    Send_IMC_Command(32'd97963751);
    Send_IMC_Command(32'd98034447);
    Send_IMC_Command(32'd299820297);
    Send_IMC_Command(32'd98700299);
    Send_IMC_Command(32'd286057230);
    Send_IMC_Command(32'd98887400);
    Send_IMC_Command(32'd300471309);
    Send_IMC_Command(32'd99083274);
    Send_IMC_Command(32'd85201536);
    Send_IMC_Command(32'd85397889);
    Send_IMC_Command(32'd85398658);
    Send_IMC_Command(32'd85398147);
    Send_IMC_Command(32'd85333397);
    Send_IMC_Command(32'd93655172);
    Send_IMC_Command(32'd92542085);
    Send_IMC_Command(32'd92373126);
    Send_IMC_Command(32'd92542855);
    Send_IMC_Command(32'd92541320);
    Send_IMC_Command(32'd92832649);
    Send_IMC_Command(32'd85165718);
    Send_IMC_Command(32'd93721226);
    Send_IMC_Command(32'd93722251);
    Send_IMC_Command(32'd92934284);
    Send_IMC_Command(32'd92968333);
    Send_IMC_Command(32'd93029006);
    Send_IMC_Command(32'd84971151);
    Send_IMC_Command(32'd93163152);
    Send_IMC_Command(32'd93160337);
    Send_IMC_Command(32'd93687442);
    Send_IMC_Command(32'd92377747);
    Send_IMC_Command(32'd85430932);
    Send_IMC_Command(32'd75926167);
    Send_IMC_Command(32'd76123288);
    Send_IMC_Command(32'd93886361);
    Send_IMC_Command(32'd75829402);
    Send_IMC_Command(32'd94017435);
    Send_IMC_Command(32'd75600540);
    Send_IMC_Command(32'd76055709);
    Send_IMC_Command(32'd94215326);
    Send_IMC_Command(32'd75992991);
    Send_IMC_Command(32'd94346400);
    Send_IMC_Command(32'd75665057);
    Send_IMC_Command(32'd75534498);
    Send_IMC_Command(32'd94544291);
    Send_IMC_Command(32'd75730340);
    Send_IMC_Command(32'd94675365);
    Send_IMC_Command(32'd93948838);
    Send_IMC_Command(32'd94086567);
    Send_IMC_Command(32'd94282664);
    Send_IMC_Command(32'd94414249);
    Send_IMC_Command(32'd94806954);
    Send_IMC_Command(32'd94867883);
    Send_IMC_Command(32'd94933932);
    Send_IMC_Command(32'd94999725);
    Send_IMC_Command(32'd95071150);
    Send_IMC_Command(32'd78294191);
    Send_IMC_Command(32'd95268784);
    Send_IMC_Command(32'd78557361);
    Send_IMC_Command(32'd95529906);
    Send_IMC_Command(32'd95202739);
    Send_IMC_Command(32'd95137716);
    Send_IMC_Command(32'd78951349);
    Send_IMC_Command(32'd95792566);
    Send_IMC_Command(32'd95205047);
    Send_IMC_Command(32'd95467192);
    Send_IMC_Command(32'd78493881);
    Send_IMC_Command(32'd96057274);
    Send_IMC_Command(32'd95467963);
    Send_IMC_Command(32'd78822332);
    Send_IMC_Command(32'd95337661);
    Send_IMC_Command(32'd96320190);
    Send_IMC_Command(32'd95598271);
    Send_IMC_Command(32'd95600064);
    Send_IMC_Command(32'd95861441);
    Send_IMC_Command(32'd96452290);
    Send_IMC_Command(32'd79792835);
    Send_IMC_Command(32'd79334596);
    Send_IMC_Command(32'd79040709);
    Send_IMC_Command(32'd79729350);
    Send_IMC_Command(32'd79529159);
    Send_IMC_Command(32'd78811080);
    Send_IMC_Command(32'd79662793);
    Send_IMC_Command(32'd79859914);
    Send_IMC_Command(32'd79597003);
    Send_IMC_Command(32'd79791820);
    Send_IMC_Command(32'd79333837);
    Send_IMC_Command(32'd79070670);
    Send_IMC_Command(32'd79725007);
    Send_IMC_Command(32'd79530192);
    Send_IMC_Command(32'd78809041);
    Send_IMC_Command(32'd79659730);
    Send_IMC_Command(32'd79855827);
    Send_IMC_Command(32'd79594452);
    Send_IMC_Command(32'd97702869);
    Send_IMC_Command(32'd97375702);
    Send_IMC_Command(32'd97310423);
    Send_IMC_Command(32'd96716248);
    Send_IMC_Command(32'd96781273);
    Send_IMC_Command(32'd96913370);
    Send_IMC_Command(32'd97507547);
    Send_IMC_Command(32'd97180380);
    Send_IMC_Command(32'd97246173);
    Send_IMC_Command(32'd98360798);
    Send_IMC_Command(32'd98228703);
    Send_IMC_Command(32'd96913632);
    Send_IMC_Command(32'd97572321);
    Send_IMC_Command(32'd98099426);
    Send_IMC_Command(32'd98033428);
    Send_IMC_Command(32'd97115363);
    Send_IMC_Command(32'd97640164);
    Send_IMC_Command(32'd98689765);
    Send_IMC_Command(32'd298837264);
    Send_IMC_Command(32'd97706982);
    Send_IMC_Command(32'd97963751);
    Send_IMC_Command(32'd98034455);
    Send_IMC_Command(32'd299820305);
    Send_IMC_Command(32'd98702355);
    Send_IMC_Command(32'd286581526);
    Send_IMC_Command(32'd98887400);
    Send_IMC_Command(32'd300471317);
    Send_IMC_Command(32'd99083282);
    Send_IMC_Command(32'd85727872);
    Send_IMC_Command(32'd85924225);
    Send_IMC_Command(32'd85924994);
    Send_IMC_Command(32'd85924483);
    Send_IMC_Command(32'd85859733);
    Send_IMC_Command(32'd93657220);
    Send_IMC_Command(32'd92544133);
    Send_IMC_Command(32'd92373126);
    Send_IMC_Command(32'd92544903);
    Send_IMC_Command(32'd92543368);
    Send_IMC_Command(32'd92832649);
    Send_IMC_Command(32'd85690006);
    Send_IMC_Command(32'd93723274);
    Send_IMC_Command(32'd93724299);
    Send_IMC_Command(32'd92936332);
    Send_IMC_Command(32'd92968333);
    Send_IMC_Command(32'd93029006);
    Send_IMC_Command(32'd85495439);
    Send_IMC_Command(32'd93163152);
    Send_IMC_Command(32'd93160337);
    Send_IMC_Command(32'd93687442);
    Send_IMC_Command(32'd92377747);
    Send_IMC_Command(32'd85955220);
    Send_IMC_Command(32'd75926167);
    Send_IMC_Command(32'd76123288);
    Send_IMC_Command(32'd93886361);
    Send_IMC_Command(32'd75831450);
    Send_IMC_Command(32'd94017435);
    Send_IMC_Command(32'd75600540);
    Send_IMC_Command(32'd76055709);
    Send_IMC_Command(32'd94215326);
    Send_IMC_Command(32'd75992991);
    Send_IMC_Command(32'd94346400);
    Send_IMC_Command(32'd75665057);
    Send_IMC_Command(32'd75534498);
    Send_IMC_Command(32'd94544291);
    Send_IMC_Command(32'd75730340);
    Send_IMC_Command(32'd94675365);
    Send_IMC_Command(32'd93948838);
    Send_IMC_Command(32'd94086567);
    Send_IMC_Command(32'd94282664);
    Send_IMC_Command(32'd94414249);
    Send_IMC_Command(32'd94806954);
    Send_IMC_Command(32'd94867883);
    Send_IMC_Command(32'd94933932);
    Send_IMC_Command(32'd94999725);
    Send_IMC_Command(32'd95071150);
    Send_IMC_Command(32'd78294191);
    Send_IMC_Command(32'd95268784);
    Send_IMC_Command(32'd78557361);
    Send_IMC_Command(32'd95529906);
    Send_IMC_Command(32'd95202739);
    Send_IMC_Command(32'd95137716);
    Send_IMC_Command(32'd78951349);
    Send_IMC_Command(32'd95792566);
    Send_IMC_Command(32'd95205047);
    Send_IMC_Command(32'd95467192);
    Send_IMC_Command(32'd78493881);
    Send_IMC_Command(32'd96057274);
    Send_IMC_Command(32'd95467963);
    Send_IMC_Command(32'd78822332);
    Send_IMC_Command(32'd95337661);
    Send_IMC_Command(32'd96320190);
    Send_IMC_Command(32'd95598271);
    Send_IMC_Command(32'd95600064);
    Send_IMC_Command(32'd95861441);
    Send_IMC_Command(32'd96452290);
    Send_IMC_Command(32'd79792835);
    Send_IMC_Command(32'd79334596);
    Send_IMC_Command(32'd79042757);
    Send_IMC_Command(32'd79729350);
    Send_IMC_Command(32'd79529159);
    Send_IMC_Command(32'd78811080);
    Send_IMC_Command(32'd79662793);
    Send_IMC_Command(32'd79859914);
    Send_IMC_Command(32'd79597003);
    Send_IMC_Command(32'd79791820);
    Send_IMC_Command(32'd79333837);
    Send_IMC_Command(32'd79070670);
    Send_IMC_Command(32'd79725007);
    Send_IMC_Command(32'd79530192);
    Send_IMC_Command(32'd78809041);
    Send_IMC_Command(32'd79659730);
    Send_IMC_Command(32'd79855827);
    Send_IMC_Command(32'd79594452);
    Send_IMC_Command(32'd97702869);
    Send_IMC_Command(32'd97375702);
    Send_IMC_Command(32'd97310423);
    Send_IMC_Command(32'd96716248);
    Send_IMC_Command(32'd96781273);
    Send_IMC_Command(32'd96913370);
    Send_IMC_Command(32'd97507547);
    Send_IMC_Command(32'd97180380);
    Send_IMC_Command(32'd97246173);
    Send_IMC_Command(32'd98360798);
    Send_IMC_Command(32'd98228703);
    Send_IMC_Command(32'd96913632);
    Send_IMC_Command(32'd97572321);
    Send_IMC_Command(32'd98099426);
    Send_IMC_Command(32'd98033436);
    Send_IMC_Command(32'd97115363);
    Send_IMC_Command(32'd97640164);
    Send_IMC_Command(32'd98689765);
    Send_IMC_Command(32'd298837272);
    Send_IMC_Command(32'd97706982);
    Send_IMC_Command(32'd97963751);
    Send_IMC_Command(32'd98034463);
    Send_IMC_Command(32'd299820313);
    Send_IMC_Command(32'd98704411);
    Send_IMC_Command(32'd287105822);
    Send_IMC_Command(32'd98887400);
    Send_IMC_Command(32'd300471325);
    Send_IMC_Command(32'd99083290);
    Send_IMC_Command(32'd86254208);
    Send_IMC_Command(32'd86450561);
    Send_IMC_Command(32'd86451330);
    Send_IMC_Command(32'd86450819);
    Send_IMC_Command(32'd86386069);
    Send_IMC_Command(32'd93659268);
    Send_IMC_Command(32'd92546181);
    Send_IMC_Command(32'd92373126);
    Send_IMC_Command(32'd92546951);
    Send_IMC_Command(32'd92545416);
    Send_IMC_Command(32'd92832649);
    Send_IMC_Command(32'd86214294);
    Send_IMC_Command(32'd93725322);
    Send_IMC_Command(32'd93726347);
    Send_IMC_Command(32'd92938380);
    Send_IMC_Command(32'd92968333);
    Send_IMC_Command(32'd93029006);
    Send_IMC_Command(32'd86019727);
    Send_IMC_Command(32'd93163152);
    Send_IMC_Command(32'd93160337);
    Send_IMC_Command(32'd93687442);
    Send_IMC_Command(32'd92377747);
    Send_IMC_Command(32'd86479508);
    Send_IMC_Command(32'd75926167);
    Send_IMC_Command(32'd76123288);
    Send_IMC_Command(32'd93886361);
    Send_IMC_Command(32'd75833498);
    Send_IMC_Command(32'd94017435);
    Send_IMC_Command(32'd75600540);
    Send_IMC_Command(32'd76055709);
    Send_IMC_Command(32'd94215326);
    Send_IMC_Command(32'd75992991);
    Send_IMC_Command(32'd94346400);
    Send_IMC_Command(32'd75665057);
    Send_IMC_Command(32'd75534498);
    Send_IMC_Command(32'd94544291);
    Send_IMC_Command(32'd75730340);
    Send_IMC_Command(32'd94675365);
    Send_IMC_Command(32'd93948838);
    Send_IMC_Command(32'd94086567);
    Send_IMC_Command(32'd94282664);
    Send_IMC_Command(32'd94414249);
    Send_IMC_Command(32'd94806954);
    Send_IMC_Command(32'd94867883);
    Send_IMC_Command(32'd94933932);
    Send_IMC_Command(32'd94999725);
    Send_IMC_Command(32'd95071150);
    Send_IMC_Command(32'd78294191);
    Send_IMC_Command(32'd95268784);
    Send_IMC_Command(32'd78557361);
    Send_IMC_Command(32'd95529906);
    Send_IMC_Command(32'd95202739);
    Send_IMC_Command(32'd95137716);
    Send_IMC_Command(32'd78951349);
    Send_IMC_Command(32'd95792566);
    Send_IMC_Command(32'd95205047);
    Send_IMC_Command(32'd95467192);
    Send_IMC_Command(32'd78493881);
    Send_IMC_Command(32'd96057274);
    Send_IMC_Command(32'd95467963);
    Send_IMC_Command(32'd78822332);
    Send_IMC_Command(32'd95337661);
    Send_IMC_Command(32'd96320190);
    Send_IMC_Command(32'd95598271);
    Send_IMC_Command(32'd95600064);
    Send_IMC_Command(32'd95861441);
    Send_IMC_Command(32'd96452290);
    Send_IMC_Command(32'd79792835);
    Send_IMC_Command(32'd79334596);
    Send_IMC_Command(32'd79044805);
    Send_IMC_Command(32'd79729350);
    Send_IMC_Command(32'd79529159);
    Send_IMC_Command(32'd78811080);
    Send_IMC_Command(32'd79662793);
    Send_IMC_Command(32'd79859914);
    Send_IMC_Command(32'd79597003);
    Send_IMC_Command(32'd79791820);
    Send_IMC_Command(32'd79333837);
    Send_IMC_Command(32'd79070670);
    Send_IMC_Command(32'd79725007);
    Send_IMC_Command(32'd79530192);
    Send_IMC_Command(32'd78809041);
    Send_IMC_Command(32'd79659730);
    Send_IMC_Command(32'd79855827);
    Send_IMC_Command(32'd79594452);
    Send_IMC_Command(32'd97702869);
    Send_IMC_Command(32'd97375702);
    Send_IMC_Command(32'd97310423);
    Send_IMC_Command(32'd96716248);
    Send_IMC_Command(32'd96781273);
    Send_IMC_Command(32'd96913370);
    Send_IMC_Command(32'd97507547);
    Send_IMC_Command(32'd97180380);
    Send_IMC_Command(32'd97246173);
    Send_IMC_Command(32'd98360798);
    Send_IMC_Command(32'd98228703);
    Send_IMC_Command(32'd96913632);
    Send_IMC_Command(32'd97572321);
    Send_IMC_Command(32'd98099426);
    Send_IMC_Command(32'd98033444);
    Send_IMC_Command(32'd97115363);
    Send_IMC_Command(32'd97640164);
    Send_IMC_Command(32'd98689765);
    Send_IMC_Command(32'd298837280);
    Send_IMC_Command(32'd97706982);
    Send_IMC_Command(32'd97963751);
    Send_IMC_Command(32'd98034471);
    Send_IMC_Command(32'd299820321);
    Send_IMC_Command(32'd98706467);
    Send_IMC_Command(32'd287630118);
    Send_IMC_Command(32'd98887400);
    Send_IMC_Command(32'd300471333);
    Send_IMC_Command(32'd99083298);
    Send_IMC_Command(32'd86780544);
    Send_IMC_Command(32'd86976897);
    Send_IMC_Command(32'd86977666);
    Send_IMC_Command(32'd86977155);
    Send_IMC_Command(32'd86912405);
    Send_IMC_Command(32'd93661316);
    Send_IMC_Command(32'd92548229);
    Send_IMC_Command(32'd92373126);
    Send_IMC_Command(32'd92548999);
    Send_IMC_Command(32'd92547464);
    Send_IMC_Command(32'd92832649);
    Send_IMC_Command(32'd86738582);
    Send_IMC_Command(32'd93727370);
    Send_IMC_Command(32'd93728395);
    Send_IMC_Command(32'd92940428);
    Send_IMC_Command(32'd92968333);
    Send_IMC_Command(32'd93029006);
    Send_IMC_Command(32'd86544015);
    Send_IMC_Command(32'd93163152);
    Send_IMC_Command(32'd93160337);
    Send_IMC_Command(32'd93687442);
    Send_IMC_Command(32'd92377747);
    Send_IMC_Command(32'd87003796);
    Send_IMC_Command(32'd75926167);
    Send_IMC_Command(32'd76123288);
    Send_IMC_Command(32'd93886361);
    Send_IMC_Command(32'd75835546);
    Send_IMC_Command(32'd94017435);
    Send_IMC_Command(32'd75600540);
    Send_IMC_Command(32'd76055709);
    Send_IMC_Command(32'd94215326);
    Send_IMC_Command(32'd75992991);
    Send_IMC_Command(32'd94346400);
    Send_IMC_Command(32'd75665057);
    Send_IMC_Command(32'd75534498);
    Send_IMC_Command(32'd94544291);
    Send_IMC_Command(32'd75730340);
    Send_IMC_Command(32'd94675365);
    Send_IMC_Command(32'd93948838);
    Send_IMC_Command(32'd94086567);
    Send_IMC_Command(32'd94282664);
    Send_IMC_Command(32'd94414249);
    Send_IMC_Command(32'd94806954);
    Send_IMC_Command(32'd94867883);
    Send_IMC_Command(32'd94933932);
    Send_IMC_Command(32'd94999725);
    Send_IMC_Command(32'd95071150);
    Send_IMC_Command(32'd78294191);
    Send_IMC_Command(32'd95268784);
    Send_IMC_Command(32'd78557361);
    Send_IMC_Command(32'd95529906);
    Send_IMC_Command(32'd95202739);
    Send_IMC_Command(32'd95137716);
    Send_IMC_Command(32'd78951349);
    Send_IMC_Command(32'd95792566);
    Send_IMC_Command(32'd95205047);
    Send_IMC_Command(32'd95467192);
    Send_IMC_Command(32'd78493881);
    Send_IMC_Command(32'd96057274);
    Send_IMC_Command(32'd95467963);
    Send_IMC_Command(32'd78822332);
    Send_IMC_Command(32'd95337661);
    Send_IMC_Command(32'd96320190);
    Send_IMC_Command(32'd95598271);
    Send_IMC_Command(32'd95600064);
    Send_IMC_Command(32'd95861441);
    Send_IMC_Command(32'd96452290);
    Send_IMC_Command(32'd79792835);
    Send_IMC_Command(32'd79334596);
    Send_IMC_Command(32'd79046853);
    Send_IMC_Command(32'd79729350);
    Send_IMC_Command(32'd79529159);
    Send_IMC_Command(32'd78811080);
    Send_IMC_Command(32'd79662793);
    Send_IMC_Command(32'd79859914);
    Send_IMC_Command(32'd79597003);
    Send_IMC_Command(32'd79791820);
    Send_IMC_Command(32'd79333837);
    Send_IMC_Command(32'd79070670);
    Send_IMC_Command(32'd79725007);
    Send_IMC_Command(32'd79530192);
    Send_IMC_Command(32'd78809041);
    Send_IMC_Command(32'd79659730);
    Send_IMC_Command(32'd79855827);
    Send_IMC_Command(32'd79594452);
    Send_IMC_Command(32'd97702869);
    Send_IMC_Command(32'd97375702);
    Send_IMC_Command(32'd97310423);
    Send_IMC_Command(32'd96716248);
    Send_IMC_Command(32'd96781273);
    Send_IMC_Command(32'd96913370);
    Send_IMC_Command(32'd97507547);
    Send_IMC_Command(32'd97180380);
    Send_IMC_Command(32'd97246173);
    Send_IMC_Command(32'd98360798);
    Send_IMC_Command(32'd98228703);
    Send_IMC_Command(32'd96913632);
    Send_IMC_Command(32'd97572321);
    Send_IMC_Command(32'd98099426);
    Send_IMC_Command(32'd98033452);
    Send_IMC_Command(32'd97115363);
    Send_IMC_Command(32'd97640164);
    Send_IMC_Command(32'd98689765);
    Send_IMC_Command(32'd298837288);
    Send_IMC_Command(32'd97706982);
    Send_IMC_Command(32'd97963751);
    Send_IMC_Command(32'd98034479);
    Send_IMC_Command(32'd299820329);
    Send_IMC_Command(32'd98708523);
    Send_IMC_Command(32'd288154414);
    Send_IMC_Command(32'd98887400);
    Send_IMC_Command(32'd300471341);
    Send_IMC_Command(32'd99083306);
    Send_IMC_Command(32'd87306880);
    Send_IMC_Command(32'd87503233);
    Send_IMC_Command(32'd87504002);
    Send_IMC_Command(32'd87503491);
    Send_IMC_Command(32'd87438741);
    Send_IMC_Command(32'd93663364);
    Send_IMC_Command(32'd92550277);
    Send_IMC_Command(32'd92373126);
    Send_IMC_Command(32'd92551047);
    Send_IMC_Command(32'd92549512);
    Send_IMC_Command(32'd92832649);
    Send_IMC_Command(32'd87262870);
    Send_IMC_Command(32'd93729418);
    Send_IMC_Command(32'd93730443);
    Send_IMC_Command(32'd92942476);
    Send_IMC_Command(32'd92968333);
    Send_IMC_Command(32'd93029006);
    Send_IMC_Command(32'd87068303);
    Send_IMC_Command(32'd93163152);
    Send_IMC_Command(32'd93160337);
    Send_IMC_Command(32'd93687442);
    Send_IMC_Command(32'd92377747);
    Send_IMC_Command(32'd87528084);
    Send_IMC_Command(32'd75926167);
    Send_IMC_Command(32'd76123288);
    Send_IMC_Command(32'd93886361);
    Send_IMC_Command(32'd75837594);
    Send_IMC_Command(32'd94017435);
    Send_IMC_Command(32'd75600540);
    Send_IMC_Command(32'd76055709);
    Send_IMC_Command(32'd94215326);
    Send_IMC_Command(32'd75992991);
    Send_IMC_Command(32'd94346400);
    Send_IMC_Command(32'd75665057);
    Send_IMC_Command(32'd75534498);
    Send_IMC_Command(32'd94544291);
    Send_IMC_Command(32'd75730340);
    Send_IMC_Command(32'd94675365);
    Send_IMC_Command(32'd93948838);
    Send_IMC_Command(32'd94086567);
    Send_IMC_Command(32'd94282664);
    Send_IMC_Command(32'd94414249);
    Send_IMC_Command(32'd94806954);
    Send_IMC_Command(32'd94867883);
    Send_IMC_Command(32'd94933932);
    Send_IMC_Command(32'd94999725);
    Send_IMC_Command(32'd95071150);
    Send_IMC_Command(32'd78294191);
    Send_IMC_Command(32'd95268784);
    Send_IMC_Command(32'd78557361);
    Send_IMC_Command(32'd95529906);
    Send_IMC_Command(32'd95202739);
    Send_IMC_Command(32'd95137716);
    Send_IMC_Command(32'd78951349);
    Send_IMC_Command(32'd95792566);
    Send_IMC_Command(32'd95205047);
    Send_IMC_Command(32'd95467192);
    Send_IMC_Command(32'd78493881);
    Send_IMC_Command(32'd96057274);
    Send_IMC_Command(32'd95467963);
    Send_IMC_Command(32'd78822332);
    Send_IMC_Command(32'd95337661);
    Send_IMC_Command(32'd96320190);
    Send_IMC_Command(32'd95598271);
    Send_IMC_Command(32'd95600064);
    Send_IMC_Command(32'd95861441);
    Send_IMC_Command(32'd96452290);
    Send_IMC_Command(32'd79792835);
    Send_IMC_Command(32'd79334596);
    Send_IMC_Command(32'd79048901);
    Send_IMC_Command(32'd79729350);
    Send_IMC_Command(32'd79529159);
    Send_IMC_Command(32'd78811080);
    Send_IMC_Command(32'd79662793);
    Send_IMC_Command(32'd79859914);
    Send_IMC_Command(32'd79597003);
    Send_IMC_Command(32'd79791820);
    Send_IMC_Command(32'd79333837);
    Send_IMC_Command(32'd79070670);
    Send_IMC_Command(32'd79725007);
    Send_IMC_Command(32'd79530192);
    Send_IMC_Command(32'd78809041);
    Send_IMC_Command(32'd79659730);
    Send_IMC_Command(32'd79855827);
    Send_IMC_Command(32'd79594452);
    Send_IMC_Command(32'd97702869);
    Send_IMC_Command(32'd97375702);
    Send_IMC_Command(32'd97310423);
    Send_IMC_Command(32'd96716248);
    Send_IMC_Command(32'd96781273);
    Send_IMC_Command(32'd96913370);
    Send_IMC_Command(32'd97507547);
    Send_IMC_Command(32'd97180380);
    Send_IMC_Command(32'd97246173);
    Send_IMC_Command(32'd98360798);
    Send_IMC_Command(32'd98228703);
    Send_IMC_Command(32'd96913632);
    Send_IMC_Command(32'd97572321);
    Send_IMC_Command(32'd98099426);
    Send_IMC_Command(32'd98033460);
    Send_IMC_Command(32'd97115363);
    Send_IMC_Command(32'd97640164);
    Send_IMC_Command(32'd98689765);
    Send_IMC_Command(32'd298837296);
    Send_IMC_Command(32'd97706982);
    Send_IMC_Command(32'd97963751);
    Send_IMC_Command(32'd98034487);
    Send_IMC_Command(32'd299820337);
    Send_IMC_Command(32'd98710579);
    Send_IMC_Command(32'd288678710);
    Send_IMC_Command(32'd98887400);
    Send_IMC_Command(32'd300471349);
    Send_IMC_Command(32'd99083314);
    Send_IMC_Command(32'd87833216);
    Send_IMC_Command(32'd88029569);
    Send_IMC_Command(32'd88030338);
    Send_IMC_Command(32'd88029827);
    Send_IMC_Command(32'd87965077);
    Send_IMC_Command(32'd93665412);
    Send_IMC_Command(32'd92552325);
    Send_IMC_Command(32'd92373126);
    Send_IMC_Command(32'd92553095);
    Send_IMC_Command(32'd92551560);
    Send_IMC_Command(32'd92832649);
    Send_IMC_Command(32'd87787158);
    Send_IMC_Command(32'd93731466);
    Send_IMC_Command(32'd93732491);
    Send_IMC_Command(32'd92944524);
    Send_IMC_Command(32'd92968333);
    Send_IMC_Command(32'd93029006);
    Send_IMC_Command(32'd87592591);
    Send_IMC_Command(32'd93163152);
    Send_IMC_Command(32'd93160337);
    Send_IMC_Command(32'd93687442);
    Send_IMC_Command(32'd92377747);
    Send_IMC_Command(32'd88052372);
    Send_IMC_Command(32'd75926167);
    Send_IMC_Command(32'd76123288);
    Send_IMC_Command(32'd93886361);
    Send_IMC_Command(32'd75839642);
    Send_IMC_Command(32'd94017435);
    Send_IMC_Command(32'd75600540);
    Send_IMC_Command(32'd76055709);
    Send_IMC_Command(32'd94215326);
    Send_IMC_Command(32'd75992991);
    Send_IMC_Command(32'd94346400);
    Send_IMC_Command(32'd75665057);
    Send_IMC_Command(32'd75534498);
    Send_IMC_Command(32'd94544291);
    Send_IMC_Command(32'd75730340);
    Send_IMC_Command(32'd94675365);
    Send_IMC_Command(32'd93948838);
    Send_IMC_Command(32'd94086567);
    Send_IMC_Command(32'd94282664);
    Send_IMC_Command(32'd94414249);
    Send_IMC_Command(32'd94806954);
    Send_IMC_Command(32'd94867883);
    Send_IMC_Command(32'd94933932);
    Send_IMC_Command(32'd94999725);
    Send_IMC_Command(32'd95071150);
    Send_IMC_Command(32'd78294191);
    Send_IMC_Command(32'd95268784);
    Send_IMC_Command(32'd78557361);
    Send_IMC_Command(32'd95529906);
    Send_IMC_Command(32'd95202739);
    Send_IMC_Command(32'd95137716);
    Send_IMC_Command(32'd78951349);
    Send_IMC_Command(32'd95792566);
    Send_IMC_Command(32'd95205047);
    Send_IMC_Command(32'd95467192);
    Send_IMC_Command(32'd78493881);
    Send_IMC_Command(32'd96057274);
    Send_IMC_Command(32'd95467963);
    Send_IMC_Command(32'd78822332);
    Send_IMC_Command(32'd95337661);
    Send_IMC_Command(32'd96320190);
    Send_IMC_Command(32'd95598271);
    Send_IMC_Command(32'd95600064);
    Send_IMC_Command(32'd95861441);
    Send_IMC_Command(32'd96452290);
    Send_IMC_Command(32'd79792835);
    Send_IMC_Command(32'd79334596);
    Send_IMC_Command(32'd79050949);
    Send_IMC_Command(32'd79729350);
    Send_IMC_Command(32'd79529159);
    Send_IMC_Command(32'd78811080);
    Send_IMC_Command(32'd79662793);
    Send_IMC_Command(32'd79859914);
    Send_IMC_Command(32'd79597003);
    Send_IMC_Command(32'd79791820);
    Send_IMC_Command(32'd79333837);
    Send_IMC_Command(32'd79070670);
    Send_IMC_Command(32'd79725007);
    Send_IMC_Command(32'd79530192);
    Send_IMC_Command(32'd78809041);
    Send_IMC_Command(32'd79659730);
    Send_IMC_Command(32'd79855827);
    Send_IMC_Command(32'd79594452);
    Send_IMC_Command(32'd97702869);
    Send_IMC_Command(32'd97375702);
    Send_IMC_Command(32'd97310423);
    Send_IMC_Command(32'd96716248);
    Send_IMC_Command(32'd96781273);
    Send_IMC_Command(32'd96913370);
    Send_IMC_Command(32'd97507547);
    Send_IMC_Command(32'd97180380);
    Send_IMC_Command(32'd97246173);
    Send_IMC_Command(32'd98360798);
    Send_IMC_Command(32'd98228703);
    Send_IMC_Command(32'd96913632);
    Send_IMC_Command(32'd97572321);
    Send_IMC_Command(32'd98099426);
    Send_IMC_Command(32'd98033468);
    Send_IMC_Command(32'd97115363);
    Send_IMC_Command(32'd97640164);
    Send_IMC_Command(32'd98689765);
    Send_IMC_Command(32'd298837304);
    Send_IMC_Command(32'd97706982);
    Send_IMC_Command(32'd97963751);
    Send_IMC_Command(32'd98034495);
    Send_IMC_Command(32'd299820345);
    Send_IMC_Command(32'd98712635);
    Send_IMC_Command(32'd289203006);
    Send_IMC_Command(32'd98887400);
    Send_IMC_Command(32'd300471357);
    Send_IMC_Command(32'd99083322);
    Send_IMC_Command(32'd88359552);
    Send_IMC_Command(32'd88555905);
    Send_IMC_Command(32'd88556674);
    Send_IMC_Command(32'd88556163);
    Send_IMC_Command(32'd88491413);
    Send_IMC_Command(32'd93667460);
    Send_IMC_Command(32'd92554373);
    Send_IMC_Command(32'd92373126);
    Send_IMC_Command(32'd92555143);
    Send_IMC_Command(32'd92553608);
    Send_IMC_Command(32'd92832649);
    Send_IMC_Command(32'd88311446);
    Send_IMC_Command(32'd93733514);
    Send_IMC_Command(32'd93734539);
    Send_IMC_Command(32'd92946572);
    Send_IMC_Command(32'd92968333);
    Send_IMC_Command(32'd93029006);
    Send_IMC_Command(32'd88116879);
    Send_IMC_Command(32'd93163152);
    Send_IMC_Command(32'd93160337);
    Send_IMC_Command(32'd93687442);
    Send_IMC_Command(32'd92377747);
    Send_IMC_Command(32'd88576660);
    Send_IMC_Command(32'd75926167);
    Send_IMC_Command(32'd76123288);
    Send_IMC_Command(32'd93886361);
    Send_IMC_Command(32'd75841690);
    Send_IMC_Command(32'd94017435);
    Send_IMC_Command(32'd75600540);
    Send_IMC_Command(32'd76055709);
    Send_IMC_Command(32'd94215326);
    Send_IMC_Command(32'd75992991);
    Send_IMC_Command(32'd94346400);
    Send_IMC_Command(32'd75665057);
    Send_IMC_Command(32'd75534498);
    Send_IMC_Command(32'd94544291);
    Send_IMC_Command(32'd75730340);
    Send_IMC_Command(32'd94675365);
    Send_IMC_Command(32'd93948838);
    Send_IMC_Command(32'd94086567);
    Send_IMC_Command(32'd94282664);
    Send_IMC_Command(32'd94414249);
    Send_IMC_Command(32'd94806954);
    Send_IMC_Command(32'd94867883);
    Send_IMC_Command(32'd94933932);
    Send_IMC_Command(32'd94999725);
    Send_IMC_Command(32'd95071150);
    Send_IMC_Command(32'd78294191);
    Send_IMC_Command(32'd95268784);
    Send_IMC_Command(32'd78557361);
    Send_IMC_Command(32'd95529906);
    Send_IMC_Command(32'd95202739);
    Send_IMC_Command(32'd95137716);
    Send_IMC_Command(32'd78951349);
    Send_IMC_Command(32'd95792566);
    Send_IMC_Command(32'd95205047);
    Send_IMC_Command(32'd95467192);
    Send_IMC_Command(32'd78493881);
    Send_IMC_Command(32'd96057274);
    Send_IMC_Command(32'd95467963);
    Send_IMC_Command(32'd78822332);
    Send_IMC_Command(32'd95337661);
    Send_IMC_Command(32'd96320190);
    Send_IMC_Command(32'd95598271);
    Send_IMC_Command(32'd95600064);
    Send_IMC_Command(32'd95861441);
    Send_IMC_Command(32'd96452290);
    Send_IMC_Command(32'd79792835);
    Send_IMC_Command(32'd79334596);
    Send_IMC_Command(32'd79052997);
    Send_IMC_Command(32'd79729350);
    Send_IMC_Command(32'd79529159);
    Send_IMC_Command(32'd78811080);
    Send_IMC_Command(32'd79662793);
    Send_IMC_Command(32'd79859914);
    Send_IMC_Command(32'd79597003);
    Send_IMC_Command(32'd79791820);
    Send_IMC_Command(32'd79333837);
    Send_IMC_Command(32'd79070670);
    Send_IMC_Command(32'd79725007);
    Send_IMC_Command(32'd79530192);
    Send_IMC_Command(32'd78809041);
    Send_IMC_Command(32'd79659730);
    Send_IMC_Command(32'd79855827);
    Send_IMC_Command(32'd79594452);
    Send_IMC_Command(32'd97702869);
    Send_IMC_Command(32'd97375702);
    Send_IMC_Command(32'd97310423);
    Send_IMC_Command(32'd96716248);
    Send_IMC_Command(32'd96781273);
    Send_IMC_Command(32'd96913370);
    Send_IMC_Command(32'd97507547);
    Send_IMC_Command(32'd97180380);
    Send_IMC_Command(32'd97246173);
    Send_IMC_Command(32'd98360798);
    Send_IMC_Command(32'd98228703);
    Send_IMC_Command(32'd96913632);
    Send_IMC_Command(32'd97572321);
    Send_IMC_Command(32'd98099426);
    Send_IMC_Command(32'd98033476);
    Send_IMC_Command(32'd97115363);
    Send_IMC_Command(32'd97640164);
    Send_IMC_Command(32'd98689765);
    Send_IMC_Command(32'd298837312);
    Send_IMC_Command(32'd97706982);
    Send_IMC_Command(32'd97963751);
    Send_IMC_Command(32'd98034503);
    Send_IMC_Command(32'd299820353);
    Send_IMC_Command(32'd98714691);
    Send_IMC_Command(32'd289727302);
    Send_IMC_Command(32'd98887400);
    Send_IMC_Command(32'd300471365);
    Send_IMC_Command(32'd99083330);
    Send_IMC_Command(32'd88885888);
    Send_IMC_Command(32'd89082241);
    Send_IMC_Command(32'd89083010);
    Send_IMC_Command(32'd89082499);
    Send_IMC_Command(32'd89017749);
    Send_IMC_Command(32'd93669508);
    Send_IMC_Command(32'd92556421);
    Send_IMC_Command(32'd92373126);
    Send_IMC_Command(32'd92557191);
    Send_IMC_Command(32'd92555656);
    Send_IMC_Command(32'd92832649);
    Send_IMC_Command(32'd88835734);
    Send_IMC_Command(32'd93735562);
    Send_IMC_Command(32'd93736587);
    Send_IMC_Command(32'd92948620);
    Send_IMC_Command(32'd92968333);
    Send_IMC_Command(32'd93029006);
    Send_IMC_Command(32'd88641167);
    Send_IMC_Command(32'd93163152);
    Send_IMC_Command(32'd93160337);
    Send_IMC_Command(32'd93687442);
    Send_IMC_Command(32'd92377747);
    Send_IMC_Command(32'd89100948);
    Send_IMC_Command(32'd75926167);
    Send_IMC_Command(32'd76123288);
    Send_IMC_Command(32'd93886361);
    Send_IMC_Command(32'd75843738);
    Send_IMC_Command(32'd94017435);
    Send_IMC_Command(32'd75600540);
    Send_IMC_Command(32'd76055709);
    Send_IMC_Command(32'd94215326);
    Send_IMC_Command(32'd75992991);
    Send_IMC_Command(32'd94346400);
    Send_IMC_Command(32'd75665057);
    Send_IMC_Command(32'd75534498);
    Send_IMC_Command(32'd94544291);
    Send_IMC_Command(32'd75730340);
    Send_IMC_Command(32'd94675365);
    Send_IMC_Command(32'd93948838);
    Send_IMC_Command(32'd94086567);
    Send_IMC_Command(32'd94282664);
    Send_IMC_Command(32'd94414249);
    Send_IMC_Command(32'd94806954);
    Send_IMC_Command(32'd94867883);
    Send_IMC_Command(32'd94933932);
    Send_IMC_Command(32'd94999725);
    Send_IMC_Command(32'd95071150);
    Send_IMC_Command(32'd78294191);
    Send_IMC_Command(32'd95268784);
    Send_IMC_Command(32'd78557361);
    Send_IMC_Command(32'd95529906);
    Send_IMC_Command(32'd95202739);
    Send_IMC_Command(32'd95137716);
    Send_IMC_Command(32'd78951349);
    Send_IMC_Command(32'd95792566);
    Send_IMC_Command(32'd95205047);
    Send_IMC_Command(32'd95467192);
    Send_IMC_Command(32'd78493881);
    Send_IMC_Command(32'd96057274);
    Send_IMC_Command(32'd95467963);
    Send_IMC_Command(32'd78822332);
    Send_IMC_Command(32'd95337661);
    Send_IMC_Command(32'd96320190);
    Send_IMC_Command(32'd95598271);
    Send_IMC_Command(32'd95600064);
    Send_IMC_Command(32'd95861441);
    Send_IMC_Command(32'd96452290);
    Send_IMC_Command(32'd79792835);
    Send_IMC_Command(32'd79334596);
    Send_IMC_Command(32'd79055045);
    Send_IMC_Command(32'd79729350);
    Send_IMC_Command(32'd79529159);
    Send_IMC_Command(32'd78811080);
    Send_IMC_Command(32'd79662793);
    Send_IMC_Command(32'd79859914);
    Send_IMC_Command(32'd79597003);
    Send_IMC_Command(32'd79791820);
    Send_IMC_Command(32'd79333837);
    Send_IMC_Command(32'd79070670);
    Send_IMC_Command(32'd79725007);
    Send_IMC_Command(32'd79530192);
    Send_IMC_Command(32'd78809041);
    Send_IMC_Command(32'd79659730);
    Send_IMC_Command(32'd79855827);
    Send_IMC_Command(32'd79594452);
    Send_IMC_Command(32'd97702869);
    Send_IMC_Command(32'd97375702);
    Send_IMC_Command(32'd97310423);
    Send_IMC_Command(32'd96716248);
    Send_IMC_Command(32'd96781273);
    Send_IMC_Command(32'd96913370);
    Send_IMC_Command(32'd97507547);
    Send_IMC_Command(32'd97180380);
    Send_IMC_Command(32'd97246173);
    Send_IMC_Command(32'd98360798);
    Send_IMC_Command(32'd98228703);
    Send_IMC_Command(32'd96913632);
    Send_IMC_Command(32'd97572321);
    Send_IMC_Command(32'd98099426);
    Send_IMC_Command(32'd98033484);
    Send_IMC_Command(32'd97115363);
    Send_IMC_Command(32'd97640164);
    Send_IMC_Command(32'd98689765);
    Send_IMC_Command(32'd298837320);
    Send_IMC_Command(32'd97706982);
    Send_IMC_Command(32'd97963751);
    Send_IMC_Command(32'd98034511);
    Send_IMC_Command(32'd299820361);
    Send_IMC_Command(32'd98716747);
    Send_IMC_Command(32'd290251598);
    Send_IMC_Command(32'd98887400);
    Send_IMC_Command(32'd300471373);
    Send_IMC_Command(32'd99083338);
    Send_IMC_Command(32'd89412224);
    Send_IMC_Command(32'd89608577);
    Send_IMC_Command(32'd89609346);
    Send_IMC_Command(32'd89608835);
    Send_IMC_Command(32'd89544085);
    Send_IMC_Command(32'd93671556);
    Send_IMC_Command(32'd92558469);
    Send_IMC_Command(32'd92373126);
    Send_IMC_Command(32'd92559239);
    Send_IMC_Command(32'd92557704);
    Send_IMC_Command(32'd92832649);
    Send_IMC_Command(32'd89360022);
    Send_IMC_Command(32'd93737610);
    Send_IMC_Command(32'd93738635);
    Send_IMC_Command(32'd92950668);
    Send_IMC_Command(32'd92968333);
    Send_IMC_Command(32'd93029006);
    Send_IMC_Command(32'd89165455);
    Send_IMC_Command(32'd93163152);
    Send_IMC_Command(32'd93160337);
    Send_IMC_Command(32'd93687442);
    Send_IMC_Command(32'd92377747);
    Send_IMC_Command(32'd89625236);
    Send_IMC_Command(32'd75926167);
    Send_IMC_Command(32'd76123288);
    Send_IMC_Command(32'd93886361);
    Send_IMC_Command(32'd75845786);
    Send_IMC_Command(32'd94017435);
    Send_IMC_Command(32'd75600540);
    Send_IMC_Command(32'd76055709);
    Send_IMC_Command(32'd94215326);
    Send_IMC_Command(32'd75992991);
    Send_IMC_Command(32'd94346400);
    Send_IMC_Command(32'd75665057);
    Send_IMC_Command(32'd75534498);
    Send_IMC_Command(32'd94544291);
    Send_IMC_Command(32'd75730340);
    Send_IMC_Command(32'd94675365);
    Send_IMC_Command(32'd93948838);
    Send_IMC_Command(32'd94086567);
    Send_IMC_Command(32'd94282664);
    Send_IMC_Command(32'd94414249);
    Send_IMC_Command(32'd94806954);
    Send_IMC_Command(32'd94867883);
    Send_IMC_Command(32'd94933932);
    Send_IMC_Command(32'd94999725);
    Send_IMC_Command(32'd95071150);
    Send_IMC_Command(32'd78294191);
    Send_IMC_Command(32'd95268784);
    Send_IMC_Command(32'd78557361);
    Send_IMC_Command(32'd95529906);
    Send_IMC_Command(32'd95202739);
    Send_IMC_Command(32'd95137716);
    Send_IMC_Command(32'd78951349);
    Send_IMC_Command(32'd95792566);
    Send_IMC_Command(32'd95205047);
    Send_IMC_Command(32'd95467192);
    Send_IMC_Command(32'd78493881);
    Send_IMC_Command(32'd96057274);
    Send_IMC_Command(32'd95467963);
    Send_IMC_Command(32'd78822332);
    Send_IMC_Command(32'd95337661);
    Send_IMC_Command(32'd96320190);
    Send_IMC_Command(32'd95598271);
    Send_IMC_Command(32'd95600064);
    Send_IMC_Command(32'd95861441);
    Send_IMC_Command(32'd96452290);
    Send_IMC_Command(32'd79792835);
    Send_IMC_Command(32'd79334596);
    Send_IMC_Command(32'd79057093);
    Send_IMC_Command(32'd79729350);
    Send_IMC_Command(32'd79529159);
    Send_IMC_Command(32'd78811080);
    Send_IMC_Command(32'd79662793);
    Send_IMC_Command(32'd79859914);
    Send_IMC_Command(32'd79597003);
    Send_IMC_Command(32'd79791820);
    Send_IMC_Command(32'd79333837);
    Send_IMC_Command(32'd79070670);
    Send_IMC_Command(32'd79725007);
    Send_IMC_Command(32'd79530192);
    Send_IMC_Command(32'd78809041);
    Send_IMC_Command(32'd79659730);
    Send_IMC_Command(32'd79855827);
    Send_IMC_Command(32'd79594452);
    Send_IMC_Command(32'd97702869);
    Send_IMC_Command(32'd97375702);
    Send_IMC_Command(32'd97310423);
    Send_IMC_Command(32'd96716248);
    Send_IMC_Command(32'd96781273);
    Send_IMC_Command(32'd96913370);
    Send_IMC_Command(32'd97507547);
    Send_IMC_Command(32'd97180380);
    Send_IMC_Command(32'd97246173);
    Send_IMC_Command(32'd98360798);
    Send_IMC_Command(32'd98228703);
    Send_IMC_Command(32'd96913632);
    Send_IMC_Command(32'd97572321);
    Send_IMC_Command(32'd98099426);
    Send_IMC_Command(32'd98033492);
    Send_IMC_Command(32'd97115363);
    Send_IMC_Command(32'd97640164);
    Send_IMC_Command(32'd98689765);
    Send_IMC_Command(32'd298837328);
    Send_IMC_Command(32'd97706982);
    Send_IMC_Command(32'd97963751);
    Send_IMC_Command(32'd98034519);
    Send_IMC_Command(32'd299820369);
    Send_IMC_Command(32'd98718803);
    Send_IMC_Command(32'd290775894);
    Send_IMC_Command(32'd98887400);
    Send_IMC_Command(32'd300471381);
    Send_IMC_Command(32'd99083346);
    Send_IMC_Command(32'd89938560);
    Send_IMC_Command(32'd90134913);
    Send_IMC_Command(32'd90135682);
    Send_IMC_Command(32'd90135171);
    Send_IMC_Command(32'd90070421);
    Send_IMC_Command(32'd93673604);
    Send_IMC_Command(32'd92560517);
    Send_IMC_Command(32'd92373126);
    Send_IMC_Command(32'd92561287);
    Send_IMC_Command(32'd92559752);
    Send_IMC_Command(32'd92832649);
    Send_IMC_Command(32'd89884310);
    Send_IMC_Command(32'd93739658);
    Send_IMC_Command(32'd93740683);
    Send_IMC_Command(32'd92952716);
    Send_IMC_Command(32'd92968333);
    Send_IMC_Command(32'd93029006);
    Send_IMC_Command(32'd89689743);
    Send_IMC_Command(32'd93163152);
    Send_IMC_Command(32'd93160337);
    Send_IMC_Command(32'd93687442);
    Send_IMC_Command(32'd92377747);
    Send_IMC_Command(32'd90149524);
    Send_IMC_Command(32'd75926167);
    Send_IMC_Command(32'd76123288);
    Send_IMC_Command(32'd93886361);
    Send_IMC_Command(32'd75847834);
    Send_IMC_Command(32'd94017435);
    Send_IMC_Command(32'd75600540);
    Send_IMC_Command(32'd76055709);
    Send_IMC_Command(32'd94215326);
    Send_IMC_Command(32'd75992991);
    Send_IMC_Command(32'd94346400);
    Send_IMC_Command(32'd75665057);
    Send_IMC_Command(32'd75534498);
    Send_IMC_Command(32'd94544291);
    Send_IMC_Command(32'd75730340);
    Send_IMC_Command(32'd94675365);
    Send_IMC_Command(32'd93948838);
    Send_IMC_Command(32'd94086567);
    Send_IMC_Command(32'd94282664);
    Send_IMC_Command(32'd94414249);
    Send_IMC_Command(32'd94806954);
    Send_IMC_Command(32'd94867883);
    Send_IMC_Command(32'd94933932);
    Send_IMC_Command(32'd94999725);
    Send_IMC_Command(32'd95071150);
    Send_IMC_Command(32'd78294191);
    Send_IMC_Command(32'd95268784);
    Send_IMC_Command(32'd78557361);
    Send_IMC_Command(32'd95529906);
    Send_IMC_Command(32'd95202739);
    Send_IMC_Command(32'd95137716);
    Send_IMC_Command(32'd78951349);
    Send_IMC_Command(32'd95792566);
    Send_IMC_Command(32'd95205047);
    Send_IMC_Command(32'd95467192);
    Send_IMC_Command(32'd78493881);
    Send_IMC_Command(32'd96057274);
    Send_IMC_Command(32'd95467963);
    Send_IMC_Command(32'd78822332);
    Send_IMC_Command(32'd95337661);
    Send_IMC_Command(32'd96320190);
    Send_IMC_Command(32'd95598271);
    Send_IMC_Command(32'd95600064);
    Send_IMC_Command(32'd95861441);
    Send_IMC_Command(32'd96452290);
    Send_IMC_Command(32'd79792835);
    Send_IMC_Command(32'd79334596);
    Send_IMC_Command(32'd79059141);
    Send_IMC_Command(32'd79729350);
    Send_IMC_Command(32'd79529159);
    Send_IMC_Command(32'd78811080);
    Send_IMC_Command(32'd79662793);
    Send_IMC_Command(32'd79859914);
    Send_IMC_Command(32'd79597003);
    Send_IMC_Command(32'd79791820);
    Send_IMC_Command(32'd79333837);
    Send_IMC_Command(32'd79070670);
    Send_IMC_Command(32'd79725007);
    Send_IMC_Command(32'd79530192);
    Send_IMC_Command(32'd78809041);
    Send_IMC_Command(32'd79659730);
    Send_IMC_Command(32'd79855827);
    Send_IMC_Command(32'd79594452);
    Send_IMC_Command(32'd97702869);
    Send_IMC_Command(32'd97375702);
    Send_IMC_Command(32'd97310423);
    Send_IMC_Command(32'd96716248);
    Send_IMC_Command(32'd96781273);
    Send_IMC_Command(32'd96913370);
    Send_IMC_Command(32'd97507547);
    Send_IMC_Command(32'd97180380);
    Send_IMC_Command(32'd97246173);
    Send_IMC_Command(32'd98360798);
    Send_IMC_Command(32'd98228703);
    Send_IMC_Command(32'd96913632);
    Send_IMC_Command(32'd97572321);
    Send_IMC_Command(32'd98099426);
    Send_IMC_Command(32'd98033500);
    Send_IMC_Command(32'd97115363);
    Send_IMC_Command(32'd97640164);
    Send_IMC_Command(32'd98689765);
    Send_IMC_Command(32'd298837336);
    Send_IMC_Command(32'd97706982);
    Send_IMC_Command(32'd97963751);
    Send_IMC_Command(32'd98034527);
    Send_IMC_Command(32'd299820377);
    Send_IMC_Command(32'd98720859);
    Send_IMC_Command(32'd291300190);
    Send_IMC_Command(32'd98887400);
    Send_IMC_Command(32'd300471389);
    Send_IMC_Command(32'd99083354);
    Send_IMC_Command(32'd90464896);
    Send_IMC_Command(32'd90661249);
    Send_IMC_Command(32'd90662018);
    Send_IMC_Command(32'd90661507);
    Send_IMC_Command(32'd90596757);
    Send_IMC_Command(32'd93675652);
    Send_IMC_Command(32'd92562565);
    Send_IMC_Command(32'd92373126);
    Send_IMC_Command(32'd92563335);
    Send_IMC_Command(32'd92561800);
    Send_IMC_Command(32'd92832649);
    Send_IMC_Command(32'd90408598);
    Send_IMC_Command(32'd93741706);
    Send_IMC_Command(32'd93742731);
    Send_IMC_Command(32'd92954764);
    Send_IMC_Command(32'd92968333);
    Send_IMC_Command(32'd93029006);
    Send_IMC_Command(32'd90214031);
    Send_IMC_Command(32'd93163152);
    Send_IMC_Command(32'd93160337);
    Send_IMC_Command(32'd93687442);
    Send_IMC_Command(32'd92377747);
    Send_IMC_Command(32'd90673812);
    Send_IMC_Command(32'd75926167);
    Send_IMC_Command(32'd76123288);
    Send_IMC_Command(32'd93886361);
    Send_IMC_Command(32'd75849882);
    Send_IMC_Command(32'd94017435);
    Send_IMC_Command(32'd75600540);
    Send_IMC_Command(32'd76055709);
    Send_IMC_Command(32'd94215326);
    Send_IMC_Command(32'd75992991);
    Send_IMC_Command(32'd94346400);
    Send_IMC_Command(32'd75665057);
    Send_IMC_Command(32'd75534498);
    Send_IMC_Command(32'd94544291);
    Send_IMC_Command(32'd75730340);
    Send_IMC_Command(32'd94675365);
    Send_IMC_Command(32'd93948838);
    Send_IMC_Command(32'd94086567);
    Send_IMC_Command(32'd94282664);
    Send_IMC_Command(32'd94414249);
    Send_IMC_Command(32'd94806954);
    Send_IMC_Command(32'd94867883);
    Send_IMC_Command(32'd94933932);
    Send_IMC_Command(32'd94999725);
    Send_IMC_Command(32'd95071150);
    Send_IMC_Command(32'd78294191);
    Send_IMC_Command(32'd95268784);
    Send_IMC_Command(32'd78557361);
    Send_IMC_Command(32'd95529906);
    Send_IMC_Command(32'd95202739);
    Send_IMC_Command(32'd95137716);
    Send_IMC_Command(32'd78951349);
    Send_IMC_Command(32'd95792566);
    Send_IMC_Command(32'd95205047);
    Send_IMC_Command(32'd95467192);
    Send_IMC_Command(32'd78493881);
    Send_IMC_Command(32'd96057274);
    Send_IMC_Command(32'd95467963);
    Send_IMC_Command(32'd78822332);
    Send_IMC_Command(32'd95337661);
    Send_IMC_Command(32'd96320190);
    Send_IMC_Command(32'd95598271);
    Send_IMC_Command(32'd95600064);
    Send_IMC_Command(32'd95861441);
    Send_IMC_Command(32'd96452290);
    Send_IMC_Command(32'd79792835);
    Send_IMC_Command(32'd79334596);
    Send_IMC_Command(32'd79061189);
    Send_IMC_Command(32'd79729350);
    Send_IMC_Command(32'd79529159);
    Send_IMC_Command(32'd78811080);
    Send_IMC_Command(32'd79662793);
    Send_IMC_Command(32'd79859914);
    Send_IMC_Command(32'd79597003);
    Send_IMC_Command(32'd79791820);
    Send_IMC_Command(32'd79333837);
    Send_IMC_Command(32'd79070670);
    Send_IMC_Command(32'd79725007);
    Send_IMC_Command(32'd79530192);
    Send_IMC_Command(32'd78809041);
    Send_IMC_Command(32'd79659730);
    Send_IMC_Command(32'd79855827);
    Send_IMC_Command(32'd79594452);
    Send_IMC_Command(32'd97702869);
    Send_IMC_Command(32'd97375702);
    Send_IMC_Command(32'd97310423);
    Send_IMC_Command(32'd96716248);
    Send_IMC_Command(32'd96781273);
    Send_IMC_Command(32'd96913370);
    Send_IMC_Command(32'd97507547);
    Send_IMC_Command(32'd97180380);
    Send_IMC_Command(32'd97246173);
    Send_IMC_Command(32'd98360798);
    Send_IMC_Command(32'd98228703);
    Send_IMC_Command(32'd96913632);
    Send_IMC_Command(32'd97572321);
    Send_IMC_Command(32'd98099426);
    Send_IMC_Command(32'd98033508);
    Send_IMC_Command(32'd97115363);
    Send_IMC_Command(32'd97640164);
    Send_IMC_Command(32'd98689765);
    Send_IMC_Command(32'd298837344);
    Send_IMC_Command(32'd97706982);
    Send_IMC_Command(32'd97963751);
    Send_IMC_Command(32'd98034535);
    Send_IMC_Command(32'd299820385);
    Send_IMC_Command(32'd98722915);
    Send_IMC_Command(32'd291824486);
    Send_IMC_Command(32'd98887400);
    Send_IMC_Command(32'd300471397);
    Send_IMC_Command(32'd99083362);
    Send_IMC_Command(32'd90991232);
    Send_IMC_Command(32'd91187585);
    Send_IMC_Command(32'd91188354);
    Send_IMC_Command(32'd91187843);
    Send_IMC_Command(32'd91123093);
    Send_IMC_Command(32'd93677700);
    Send_IMC_Command(32'd92564613);
    Send_IMC_Command(32'd92373126);
    Send_IMC_Command(32'd92565383);
    Send_IMC_Command(32'd92563848);
    Send_IMC_Command(32'd92832649);
    Send_IMC_Command(32'd90932886);
    Send_IMC_Command(32'd93743754);
    Send_IMC_Command(32'd93744779);
    Send_IMC_Command(32'd92956812);
    Send_IMC_Command(32'd92968333);
    Send_IMC_Command(32'd93029006);
    Send_IMC_Command(32'd90738319);
    Send_IMC_Command(32'd93163152);
    Send_IMC_Command(32'd93160337);
    Send_IMC_Command(32'd93687442);
    Send_IMC_Command(32'd92377747);
    Send_IMC_Command(32'd91198100);
    Send_IMC_Command(32'd75926167);
    Send_IMC_Command(32'd76123288);
    Send_IMC_Command(32'd93886361);
    Send_IMC_Command(32'd75851930);
    Send_IMC_Command(32'd94017435);
    Send_IMC_Command(32'd75600540);
    Send_IMC_Command(32'd76055709);
    Send_IMC_Command(32'd94215326);
    Send_IMC_Command(32'd75992991);
    Send_IMC_Command(32'd94346400);
    Send_IMC_Command(32'd75665057);
    Send_IMC_Command(32'd75534498);
    Send_IMC_Command(32'd94544291);
    Send_IMC_Command(32'd75730340);
    Send_IMC_Command(32'd94675365);
    Send_IMC_Command(32'd93948838);
    Send_IMC_Command(32'd94086567);
    Send_IMC_Command(32'd94282664);
    Send_IMC_Command(32'd94414249);
    Send_IMC_Command(32'd94806954);
    Send_IMC_Command(32'd94867883);
    Send_IMC_Command(32'd94933932);
    Send_IMC_Command(32'd94999725);
    Send_IMC_Command(32'd95071150);
    Send_IMC_Command(32'd78294191);
    Send_IMC_Command(32'd95268784);
    Send_IMC_Command(32'd78557361);
    Send_IMC_Command(32'd95529906);
    Send_IMC_Command(32'd95202739);
    Send_IMC_Command(32'd95137716);
    Send_IMC_Command(32'd78951349);
    Send_IMC_Command(32'd95792566);
    Send_IMC_Command(32'd95205047);
    Send_IMC_Command(32'd95467192);
    Send_IMC_Command(32'd78493881);
    Send_IMC_Command(32'd96057274);
    Send_IMC_Command(32'd95467963);
    Send_IMC_Command(32'd78822332);
    Send_IMC_Command(32'd95337661);
    Send_IMC_Command(32'd96320190);
    Send_IMC_Command(32'd95598271);
    Send_IMC_Command(32'd95600064);
    Send_IMC_Command(32'd95861441);
    Send_IMC_Command(32'd96452290);
    Send_IMC_Command(32'd79792835);
    Send_IMC_Command(32'd79334596);
    Send_IMC_Command(32'd79063237);
    Send_IMC_Command(32'd79729350);
    Send_IMC_Command(32'd79529159);
    Send_IMC_Command(32'd78811080);
    Send_IMC_Command(32'd79662793);
    Send_IMC_Command(32'd79859914);
    Send_IMC_Command(32'd79597003);
    Send_IMC_Command(32'd79791820);
    Send_IMC_Command(32'd79333837);
    Send_IMC_Command(32'd79070670);
    Send_IMC_Command(32'd79725007);
    Send_IMC_Command(32'd79530192);
    Send_IMC_Command(32'd78809041);
    Send_IMC_Command(32'd79659730);
    Send_IMC_Command(32'd79855827);
    Send_IMC_Command(32'd79594452);
    Send_IMC_Command(32'd97702869);
    Send_IMC_Command(32'd97375702);
    Send_IMC_Command(32'd97310423);
    Send_IMC_Command(32'd96716248);
    Send_IMC_Command(32'd96781273);
    Send_IMC_Command(32'd96913370);
    Send_IMC_Command(32'd97507547);
    Send_IMC_Command(32'd97180380);
    Send_IMC_Command(32'd97246173);
    Send_IMC_Command(32'd98360798);
    Send_IMC_Command(32'd98228703);
    Send_IMC_Command(32'd96913632);
    Send_IMC_Command(32'd97572321);
    Send_IMC_Command(32'd98099426);
    Send_IMC_Command(32'd98033516);
    Send_IMC_Command(32'd97115363);
    Send_IMC_Command(32'd97640164);
    Send_IMC_Command(32'd98689765);
    Send_IMC_Command(32'd298837352);
    Send_IMC_Command(32'd97706982);
    Send_IMC_Command(32'd97963751);
    Send_IMC_Command(32'd98034543);
    Send_IMC_Command(32'd299820393);
    Send_IMC_Command(32'd98724971);
    Send_IMC_Command(32'd292348782);
    Send_IMC_Command(32'd98887400);
    Send_IMC_Command(32'd300471405);
    Send_IMC_Command(32'd99083370);
    Send_IMC_Command(32'd91517568);
    Send_IMC_Command(32'd91713921);
    Send_IMC_Command(32'd91714690);
    Send_IMC_Command(32'd91714179);
    Send_IMC_Command(32'd91649429);
    Send_IMC_Command(32'd93679748);
    Send_IMC_Command(32'd92566661);
    Send_IMC_Command(32'd92373126);
    Send_IMC_Command(32'd92567431);
    Send_IMC_Command(32'd92565896);
    Send_IMC_Command(32'd92832649);
    Send_IMC_Command(32'd91457174);
    Send_IMC_Command(32'd93745802);
    Send_IMC_Command(32'd93746827);
    Send_IMC_Command(32'd92958860);
    Send_IMC_Command(32'd92968333);
    Send_IMC_Command(32'd93029006);
    Send_IMC_Command(32'd91262607);
    Send_IMC_Command(32'd93163152);
    Send_IMC_Command(32'd93160337);
    Send_IMC_Command(32'd93687442);
    Send_IMC_Command(32'd92377747);
    Send_IMC_Command(32'd91722388);
    Send_IMC_Command(32'd75926167);
    Send_IMC_Command(32'd76123288);
    Send_IMC_Command(32'd93886361);
    Send_IMC_Command(32'd75853978);
    Send_IMC_Command(32'd94017435);
    Send_IMC_Command(32'd75600540);
    Send_IMC_Command(32'd76055709);
    Send_IMC_Command(32'd94215326);
    Send_IMC_Command(32'd75992991);
    Send_IMC_Command(32'd94346400);
    Send_IMC_Command(32'd75665057);
    Send_IMC_Command(32'd75534498);
    Send_IMC_Command(32'd94544291);
    Send_IMC_Command(32'd75730340);
    Send_IMC_Command(32'd94675365);
    Send_IMC_Command(32'd93948838);
    Send_IMC_Command(32'd94086567);
    Send_IMC_Command(32'd94282664);
    Send_IMC_Command(32'd94414249);
    Send_IMC_Command(32'd94806954);
    Send_IMC_Command(32'd94867883);
    Send_IMC_Command(32'd94933932);
    Send_IMC_Command(32'd94999725);
    Send_IMC_Command(32'd95071150);
    Send_IMC_Command(32'd78294191);
    Send_IMC_Command(32'd95268784);
    Send_IMC_Command(32'd78557361);
    Send_IMC_Command(32'd95529906);
    Send_IMC_Command(32'd95202739);
    Send_IMC_Command(32'd95137716);
    Send_IMC_Command(32'd78951349);
    Send_IMC_Command(32'd95792566);
    Send_IMC_Command(32'd95205047);
    Send_IMC_Command(32'd95467192);
    Send_IMC_Command(32'd78493881);
    Send_IMC_Command(32'd96057274);
    Send_IMC_Command(32'd95467963);
    Send_IMC_Command(32'd78822332);
    Send_IMC_Command(32'd95337661);
    Send_IMC_Command(32'd96320190);
    Send_IMC_Command(32'd95598271);
    Send_IMC_Command(32'd95600064);
    Send_IMC_Command(32'd95861441);
    Send_IMC_Command(32'd96452290);
    Send_IMC_Command(32'd79792835);
    Send_IMC_Command(32'd79334596);
    Send_IMC_Command(32'd79065285);
    Send_IMC_Command(32'd79729350);
    Send_IMC_Command(32'd79529159);
    Send_IMC_Command(32'd78811080);
    Send_IMC_Command(32'd79662793);
    Send_IMC_Command(32'd79859914);
    Send_IMC_Command(32'd79597003);
    Send_IMC_Command(32'd79791820);
    Send_IMC_Command(32'd79333837);
    Send_IMC_Command(32'd79070670);
    Send_IMC_Command(32'd79725007);
    Send_IMC_Command(32'd79530192);
    Send_IMC_Command(32'd78809041);
    Send_IMC_Command(32'd79659730);
    Send_IMC_Command(32'd79855827);
    Send_IMC_Command(32'd79594452);
    Send_IMC_Command(32'd97702869);
    Send_IMC_Command(32'd97375702);
    Send_IMC_Command(32'd97310423);
    Send_IMC_Command(32'd96716248);
    Send_IMC_Command(32'd96781273);
    Send_IMC_Command(32'd96913370);
    Send_IMC_Command(32'd97507547);
    Send_IMC_Command(32'd97180380);
    Send_IMC_Command(32'd97246173);
    Send_IMC_Command(32'd98360798);
    Send_IMC_Command(32'd98228703);
    Send_IMC_Command(32'd96913632);
    Send_IMC_Command(32'd97572321);
    Send_IMC_Command(32'd98099426);
    Send_IMC_Command(32'd98033524);
    Send_IMC_Command(32'd97115363);
    Send_IMC_Command(32'd97640164);
    Send_IMC_Command(32'd98689765);
    Send_IMC_Command(32'd298837360);
    Send_IMC_Command(32'd97706982);
    Send_IMC_Command(32'd97963751);
    Send_IMC_Command(32'd98034551);
    Send_IMC_Command(32'd299820401);
    Send_IMC_Command(32'd98727027);
    Send_IMC_Command(32'd292873078);
    Send_IMC_Command(32'd98887400);
    Send_IMC_Command(32'd300471413);
    Send_IMC_Command(32'd99083378);
    Send_IMC_Command(32'd92043904);
    Send_IMC_Command(32'd92240257);
    Send_IMC_Command(32'd92241026);
    Send_IMC_Command(32'd92240515);
    Send_IMC_Command(32'd92175765);
    Send_IMC_Command(32'd93681796);
    Send_IMC_Command(32'd92568709);
    Send_IMC_Command(32'd92373126);
    Send_IMC_Command(32'd92569479);
    Send_IMC_Command(32'd92567944);
    Send_IMC_Command(32'd92832649);
    Send_IMC_Command(32'd91981462);
    Send_IMC_Command(32'd93747850);
    Send_IMC_Command(32'd93748875);
    Send_IMC_Command(32'd92960908);
    Send_IMC_Command(32'd92968333);
    Send_IMC_Command(32'd93029006);
    Send_IMC_Command(32'd91786895);
    Send_IMC_Command(32'd93163152);
    Send_IMC_Command(32'd93160337);
    Send_IMC_Command(32'd93687442);
    Send_IMC_Command(32'd92377747);
    Send_IMC_Command(32'd92246676);
    Send_IMC_Command(32'd75926167);
    Send_IMC_Command(32'd76123288);
    Send_IMC_Command(32'd93886361);
    Send_IMC_Command(32'd75856026);
    Send_IMC_Command(32'd94017435);
    Send_IMC_Command(32'd75600540);
    Send_IMC_Command(32'd76055709);
    Send_IMC_Command(32'd94215326);
    Send_IMC_Command(32'd75992991);
    Send_IMC_Command(32'd94346400);
    Send_IMC_Command(32'd75665057);
    Send_IMC_Command(32'd75534498);
    Send_IMC_Command(32'd94544291);
    Send_IMC_Command(32'd75730340);
    Send_IMC_Command(32'd94675365);
    Send_IMC_Command(32'd93948838);
    Send_IMC_Command(32'd94086567);
    Send_IMC_Command(32'd94282664);
    Send_IMC_Command(32'd94414249);
    Send_IMC_Command(32'd94806954);
    Send_IMC_Command(32'd94867883);
    Send_IMC_Command(32'd94933932);
    Send_IMC_Command(32'd94999725);
    Send_IMC_Command(32'd95071150);
    Send_IMC_Command(32'd78294191);
    Send_IMC_Command(32'd95268784);
    Send_IMC_Command(32'd78557361);
    Send_IMC_Command(32'd95529906);
    Send_IMC_Command(32'd95202739);
    Send_IMC_Command(32'd95137716);
    Send_IMC_Command(32'd78951349);
    Send_IMC_Command(32'd95792566);
    Send_IMC_Command(32'd95205047);
    Send_IMC_Command(32'd95467192);
    Send_IMC_Command(32'd78493881);
    Send_IMC_Command(32'd96057274);
    Send_IMC_Command(32'd95467963);
    Send_IMC_Command(32'd78822332);
    Send_IMC_Command(32'd95337661);
    Send_IMC_Command(32'd96320190);
    Send_IMC_Command(32'd95598271);
    Send_IMC_Command(32'd95600064);
    Send_IMC_Command(32'd95861441);
    Send_IMC_Command(32'd96452290);
    Send_IMC_Command(32'd79792835);
    Send_IMC_Command(32'd79334596);
    Send_IMC_Command(32'd79067333);
    Send_IMC_Command(32'd79729350);
    Send_IMC_Command(32'd79529159);
    Send_IMC_Command(32'd78811080);
    Send_IMC_Command(32'd79662793);
    Send_IMC_Command(32'd79859914);
    Send_IMC_Command(32'd79597003);
    Send_IMC_Command(32'd79791820);
    Send_IMC_Command(32'd79333837);
    Send_IMC_Command(32'd79070670);
    Send_IMC_Command(32'd79725007);
    Send_IMC_Command(32'd79530192);
    Send_IMC_Command(32'd78809041);
    Send_IMC_Command(32'd79659730);
    Send_IMC_Command(32'd79855827);
    Send_IMC_Command(32'd79594452);
    Send_IMC_Command(32'd97702869);
    Send_IMC_Command(32'd97375702);
    Send_IMC_Command(32'd97310423);
    Send_IMC_Command(32'd96716248);
    Send_IMC_Command(32'd96781273);
    Send_IMC_Command(32'd96913370);
    Send_IMC_Command(32'd97507547);
    Send_IMC_Command(32'd97180380);
    Send_IMC_Command(32'd97246173);
    Send_IMC_Command(32'd98360798);
    Send_IMC_Command(32'd98228703);
    Send_IMC_Command(32'd96913632);
    Send_IMC_Command(32'd97572321);
    Send_IMC_Command(32'd98099426);
    Send_IMC_Command(32'd98033532);
    Send_IMC_Command(32'd97115363);
    Send_IMC_Command(32'd97640164);
    Send_IMC_Command(32'd98689765);
    Send_IMC_Command(32'd298837368);
    Send_IMC_Command(32'd97706982);
    Send_IMC_Command(32'd97963751);
    Send_IMC_Command(32'd98034559);
    Send_IMC_Command(32'd299820409);
    Send_IMC_Command(32'd98729083);
    Send_IMC_Command(32'd293397374);
    Send_IMC_Command(32'd98887400);
    Send_IMC_Command(32'd300471421);
    Send_IMC_Command(32'd99083386);
endtask

task AES_MC();

    Send_IMC_Command(32'd83896480);
    Send_IMC_Command(32'd89159841);
    Send_IMC_Command(32'd83962274);
    Send_IMC_Command(32'd89225635);
    Send_IMC_Command(32'd84028068);
    Send_IMC_Command(32'd89291429);
    Send_IMC_Command(32'd84093862);
    Send_IMC_Command(32'd89357223);
    Send_IMC_Command(32'd84159656);
    Send_IMC_Command(32'd89423017);
    Send_IMC_Command(32'd84225450);
    Send_IMC_Command(32'd89488811);
    Send_IMC_Command(32'd84291244);
    Send_IMC_Command(32'd89554605);
    Send_IMC_Command(32'd89620398);
    Send_IMC_Command(32'd84357039);
    Send_IMC_Command(32'd86548912);
    Send_IMC_Command(32'd95400064);
    Send_IMC_Command(32'd84367281);
    Send_IMC_Command(32'd91791538);
    Send_IMC_Command(32'd95335056);
    Send_IMC_Command(32'd94474419);
    Send_IMC_Command(32'd95531928);
    Send_IMC_Command(32'd91991732);
    Send_IMC_Command(32'd94404789);
    Send_IMC_Command(32'd95532424);
    Send_IMC_Command(32'd94745782);
    Send_IMC_Command(32'd94811795);
    Send_IMC_Command(32'd86749111);
    Send_IMC_Command(32'd94877624);
    Send_IMC_Command(32'd94681219);
    Send_IMC_Command(32'd84038329);
    Send_IMC_Command(32'd95533498);
    Send_IMC_Command(32'd95008699);
    Send_IMC_Command(32'd94942396);
    Send_IMC_Command(32'd86680253);
    Send_IMC_Command(32'd94748034);
    Send_IMC_Command(32'd91923390);
    Send_IMC_Command(32'd94682770);
    Send_IMC_Command(32'd86604223);
    Send_IMC_Command(32'd96059328);
    Send_IMC_Command(32'd96387210);
    Send_IMC_Command(32'd96321690);
    Send_IMC_Command(32'd83997377);
    Send_IMC_Command(32'd92187586);
    Send_IMC_Command(32'd95208086);
    Send_IMC_Command(32'd86945219);
    Send_IMC_Command(32'd95077254);
    Send_IMC_Command(32'd84235716);
    Send_IMC_Command(32'd92189125);
    Send_IMC_Command(32'd89239750);
    Send_IMC_Command(32'd86878407);
    Send_IMC_Command(32'd95143813);
    Send_IMC_Command(32'd86820040);
    Send_IMC_Command(32'd92121545);
    Send_IMC_Command(32'd95078805);
    Send_IMC_Command(32'd92063946);
    Send_IMC_Command(32'd97110669);
    Send_IMC_Command(32'd96979613);
    Send_IMC_Command(32'd87010507);
    Send_IMC_Command(32'd95341447);
    Send_IMC_Command(32'd86951372);
    Send_IMC_Command(32'd97242271);
    Send_IMC_Command(32'd92253645);
    Send_IMC_Command(32'd97308047);
    Send_IMC_Command(32'd95407511);
    Send_IMC_Command(32'd95208654);
    Send_IMC_Command(32'd92720782);
    Send_IMC_Command(32'd96453071);
    Send_IMC_Command(32'd95670161);
    Send_IMC_Command(32'd94798800);
    Send_IMC_Command(32'd96129163);
    Send_IMC_Command(32'd94553809);
    Send_IMC_Command(32'd93901209);
    Send_IMC_Command(32'd94868434);
    Send_IMC_Command(32'd96129691);
    Send_IMC_Command(32'd89575123);
    Send_IMC_Command(32'd95146910);
    Send_IMC_Command(32'd89373908);
    Send_IMC_Command(32'd92066964);
    Send_IMC_Command(32'd84130773);
    Send_IMC_Command(32'd86824324);
    Send_IMC_Command(32'd94618070);
    Send_IMC_Command(32'd92853897);
    Send_IMC_Command(32'd95797207);
    Send_IMC_Command(32'd96917377);
    Send_IMC_Command(32'd84193752);
    Send_IMC_Command(32'd89381081);
    Send_IMC_Command(32'd96197004);
    Send_IMC_Command(32'd84131034);
    Send_IMC_Command(32'd95541979);
    Send_IMC_Command(32'd89447324);
    Send_IMC_Command(32'd86001856);
    Send_IMC_Command(32'd91232449);
    Send_IMC_Command(32'd86067650);
    Send_IMC_Command(32'd91298243);
    Send_IMC_Command(32'd86133444);
    Send_IMC_Command(32'd91364037);
    Send_IMC_Command(32'd86199238);
    Send_IMC_Command(32'd91429831);
    Send_IMC_Command(32'd86265032);
    Send_IMC_Command(32'd91495625);
    Send_IMC_Command(32'd86330826);
    Send_IMC_Command(32'd91561419);
    Send_IMC_Command(32'd86396620);
    Send_IMC_Command(32'd91627213);
    Send_IMC_Command(32'd91693006);
    Send_IMC_Command(32'd86462415);
    Send_IMC_Command(32'd88654288);
    Send_IMC_Command(32'd97505440);
    Send_IMC_Command(32'd86472657);
    Send_IMC_Command(32'd85508306);
    Send_IMC_Command(32'd97440432);
    Send_IMC_Command(32'd96579795);
    Send_IMC_Command(32'd97637304);
    Send_IMC_Command(32'd85708500);
    Send_IMC_Command(32'd96510165);
    Send_IMC_Command(32'd97637800);
    Send_IMC_Command(32'd96851158);
    Send_IMC_Command(32'd96917171);
    Send_IMC_Command(32'd88854487);
    Send_IMC_Command(32'd96983000);
    Send_IMC_Command(32'd96786595);
    Send_IMC_Command(32'd86143705);
    Send_IMC_Command(32'd97638874);
    Send_IMC_Command(32'd97114075);
    Send_IMC_Command(32'd97047772);
    Send_IMC_Command(32'd88785629);
    Send_IMC_Command(32'd96853410);
    Send_IMC_Command(32'd85640158);
    Send_IMC_Command(32'd96788146);
    Send_IMC_Command(32'd88676831);
    Send_IMC_Command(32'd98164704);
    Send_IMC_Command(32'd98492586);
    Send_IMC_Command(32'd98427066);
    Send_IMC_Command(32'd86102753);
    Send_IMC_Command(32'd85904354);
    Send_IMC_Command(32'd97313462);
    Send_IMC_Command(32'd89050595);
    Send_IMC_Command(32'd97182630);
    Send_IMC_Command(32'd86341092);
    Send_IMC_Command(32'd85905893);
    Send_IMC_Command(32'd91345126);
    Send_IMC_Command(32'd88983783);
    Send_IMC_Command(32'd97249189);
    Send_IMC_Command(32'd88925416);
    Send_IMC_Command(32'd85838313);
    Send_IMC_Command(32'd97184181);
    Send_IMC_Command(32'd85780714);
    Send_IMC_Command(32'd99216045);
    Send_IMC_Command(32'd99084989);
    Send_IMC_Command(32'd89115883);
    Send_IMC_Command(32'd97446823);
    Send_IMC_Command(32'd89056748);
    Send_IMC_Command(32'd99347647);
    Send_IMC_Command(32'd85970413);
    Send_IMC_Command(32'd99413423);
    Send_IMC_Command(32'd97512887);
    Send_IMC_Command(32'd97314030);
    Send_IMC_Command(32'd94826158);
    Send_IMC_Command(32'd98558447);
    Send_IMC_Command(32'd97775537);
    Send_IMC_Command(32'd96904176);
    Send_IMC_Command(32'd98234539);
    Send_IMC_Command(32'd96659185);
    Send_IMC_Command(32'd96006585);
    Send_IMC_Command(32'd96973810);
    Send_IMC_Command(32'd98235067);
    Send_IMC_Command(32'd91680499);
    Send_IMC_Command(32'd97252286);
    Send_IMC_Command(32'd91479284);
    Send_IMC_Command(32'd85783732);
    Send_IMC_Command(32'd86236149);
    Send_IMC_Command(32'd88929700);
    Send_IMC_Command(32'd96723446);
    Send_IMC_Command(32'd94959273);
    Send_IMC_Command(32'd97902583);
    Send_IMC_Command(32'd99022753);
    Send_IMC_Command(32'd86299128);
    Send_IMC_Command(32'd91486457);
    Send_IMC_Command(32'd98302380);
    Send_IMC_Command(32'd86236410);
    Send_IMC_Command(32'd97647355);
    Send_IMC_Command(32'd91552700);
    Send_IMC_Command(32'd88107232);
    Send_IMC_Command(32'd84949217);
    Send_IMC_Command(32'd88173026);
    Send_IMC_Command(32'd85015011);
    Send_IMC_Command(32'd88238820);
    Send_IMC_Command(32'd85080805);
    Send_IMC_Command(32'd88304614);
    Send_IMC_Command(32'd85146599);
    Send_IMC_Command(32'd88370408);
    Send_IMC_Command(32'd85212393);
    Send_IMC_Command(32'd88436202);
    Send_IMC_Command(32'd85278187);
    Send_IMC_Command(32'd88501996);
    Send_IMC_Command(32'd85343981);
    Send_IMC_Command(32'd85409774);
    Send_IMC_Command(32'd88567791);
    Send_IMC_Command(32'd90759664);
    Send_IMC_Command(32'd99610816);
    Send_IMC_Command(32'd88545265);
    Send_IMC_Command(32'd87613682);
    Send_IMC_Command(32'd99545808);
    Send_IMC_Command(32'd98685171);
    Send_IMC_Command(32'd99742680);
    Send_IMC_Command(32'd87813876);
    Send_IMC_Command(32'd98615541);
    Send_IMC_Command(32'd99743176);
    Send_IMC_Command(32'd98956534);
    Send_IMC_Command(32'd99022547);
    Send_IMC_Command(32'd90959863);
    Send_IMC_Command(32'd99088376);
    Send_IMC_Command(32'd98891971);
    Send_IMC_Command(32'd88216313);
    Send_IMC_Command(32'd99744250);
    Send_IMC_Command(32'd99219451);
    Send_IMC_Command(32'd99153148);
    Send_IMC_Command(32'd90891005);
    Send_IMC_Command(32'd98958786);
    Send_IMC_Command(32'd87745534);
    Send_IMC_Command(32'd98893522);
    Send_IMC_Command(32'd90782207);
    Send_IMC_Command(32'd100269824);
    Send_IMC_Command(32'd100532426);
    Send_IMC_Command(32'd100466906);
    Send_IMC_Command(32'd88207873);
    Send_IMC_Command(32'd88009474);
    Send_IMC_Command(32'd99353302);
    Send_IMC_Command(32'd91155715);
    Send_IMC_Command(32'd99222470);
    Send_IMC_Command(32'd88413444);
    Send_IMC_Command(32'd88011013);
    Send_IMC_Command(32'd85061638);
    Send_IMC_Command(32'd91088903);
    Send_IMC_Command(32'd99289029);
    Send_IMC_Command(32'd90965032);
    Send_IMC_Command(32'd87943465);
    Send_IMC_Command(32'd99232213);
    Send_IMC_Command(32'd87828522);
    Send_IMC_Command(32'd86584013);
    Send_IMC_Command(32'd84355805);
    Send_IMC_Command(32'd91221035);
    Send_IMC_Command(32'd99494855);
    Send_IMC_Command(32'd91096364);
    Send_IMC_Command(32'd86715615);
    Send_IMC_Command(32'd88075565);
    Send_IMC_Command(32'd86781391);
    Send_IMC_Command(32'd99560919);
    Send_IMC_Command(32'd99353646);
    Send_IMC_Command(32'd96874190);
    Send_IMC_Command(32'd100598063);
    Send_IMC_Command(32'd99823569);
    Send_IMC_Command(32'd99009360);
    Send_IMC_Command(32'd100290763);
    Send_IMC_Command(32'd98698833);
    Send_IMC_Command(32'd98062809);
    Send_IMC_Command(32'd99078994);
    Send_IMC_Command(32'd100291291);
    Send_IMC_Command(32'd85339731);
    Send_IMC_Command(32'd99308510);
    Send_IMC_Command(32'd85195860);
    Send_IMC_Command(32'd87839956);
    Send_IMC_Command(32'd88341333);
    Send_IMC_Command(32'd90985924);
    Send_IMC_Command(32'd98763094);
    Send_IMC_Command(32'd97015497);
    Send_IMC_Command(32'd100007767);
    Send_IMC_Command(32'd84301761);
    Send_IMC_Command(32'd88404344);
    Send_IMC_Command(32'd85162105);
    Send_IMC_Command(32'd100366796);
    Send_IMC_Command(32'd88341626);
    Send_IMC_Command(32'd99711611);
    Send_IMC_Command(32'd85228508);
    Send_IMC_Command(32'd90179584);
    Send_IMC_Command(32'd87054337);
    Send_IMC_Command(32'd90245378);
    Send_IMC_Command(32'd87120131);
    Send_IMC_Command(32'd90311172);
    Send_IMC_Command(32'd87185925);
    Send_IMC_Command(32'd90376966);
    Send_IMC_Command(32'd87251719);
    Send_IMC_Command(32'd90442792);
    Send_IMC_Command(32'd87317545);
    Send_IMC_Command(32'd90508586);
    Send_IMC_Command(32'd87383339);
    Send_IMC_Command(32'd90574380);
    Send_IMC_Command(32'd87449133);
    Send_IMC_Command(32'd87514926);
    Send_IMC_Command(32'd90640175);
    Send_IMC_Command(32'd84410704);
    Send_IMC_Command(32'd86986976);
    Send_IMC_Command(32'd90650449);
    Send_IMC_Command(32'd89653330);
    Send_IMC_Command(32'd86921968);
    Send_IMC_Command(32'd84013139);
    Send_IMC_Command(32'd89215992);
    Send_IMC_Command(32'd89861716);
    Send_IMC_Command(32'd83943509);
    Send_IMC_Command(32'd89216488);
    Send_IMC_Command(32'd84235350);
    Send_IMC_Command(32'd84301555);
    Send_IMC_Command(32'd84619095);
    Send_IMC_Command(32'd84367224);
    Send_IMC_Command(32'd84179171);
    Send_IMC_Command(32'd90321529);
    Send_IMC_Command(32'd89225594);
    Send_IMC_Command(32'd86595451);
    Send_IMC_Command(32'd86529148);
    Send_IMC_Command(32'd84542077);
    Send_IMC_Command(32'd84245986);
    Send_IMC_Command(32'd89785214);
    Send_IMC_Command(32'd84180722);
    Send_IMC_Command(32'd84498815);
    Send_IMC_Command(32'd91848480);
    Send_IMC_Command(32'd92152042);
    Send_IMC_Command(32'd92086522);
    Send_IMC_Command(32'd90264097);
    Send_IMC_Command(32'd90057506);
    Send_IMC_Command(32'd86778614);
    Send_IMC_Command(32'd84815139);
    Send_IMC_Command(32'd86647782);
    Send_IMC_Command(32'd90518820);
    Send_IMC_Command(32'd90067237);
    Send_IMC_Command(32'd87117862);
    Send_IMC_Command(32'd84748327);
    Send_IMC_Command(32'd86714341);
    Send_IMC_Command(32'd84681800);
    Send_IMC_Command(32'd89991497);
    Send_IMC_Command(32'd86657525);
    Send_IMC_Command(32'd89933898);
    Send_IMC_Command(32'd88689389);
    Send_IMC_Command(32'd86461181);
    Send_IMC_Command(32'd84880459);
    Send_IMC_Command(32'd86920167);
    Send_IMC_Command(32'd84813132);
    Send_IMC_Command(32'd88820991);
    Send_IMC_Command(32'd90123597);
    Send_IMC_Command(32'd88886767);
    Send_IMC_Command(32'd86986231);
    Send_IMC_Command(32'd86778958);
    Send_IMC_Command(32'd98979566);
    Send_IMC_Command(32'd92217679);
    Send_IMC_Command(32'd89346033);
    Send_IMC_Command(32'd84337520);
    Send_IMC_Command(32'd91910379);
    Send_IMC_Command(32'd84026993);
    Send_IMC_Command(32'd100168185);
    Send_IMC_Command(32'd84407154);
    Send_IMC_Command(32'd91910907);
    Send_IMC_Command(32'd87445107);
    Send_IMC_Command(32'd86733822);
    Send_IMC_Command(32'd87260276);
    Send_IMC_Command(32'd89945332);
    Send_IMC_Command(32'd90405749);
    Send_IMC_Command(32'd84702692);
    Send_IMC_Command(32'd84091254);
    Send_IMC_Command(32'd99120873);
    Send_IMC_Command(32'd89489271);
    Send_IMC_Command(32'd86407137);
    Send_IMC_Command(32'd90460440);
    Send_IMC_Command(32'd87234585);
    Send_IMC_Command(32'd91953644);
    Send_IMC_Command(32'd90405914);
    Send_IMC_Command(32'd89201179);
    Send_IMC_Command(32'd87301116);

endtask

task AES_Inv_SBOX();

    Send_IMC_Command(32'd92767232);
    Send_IMC_Command(32'd294028289);
    Send_IMC_Command(32'd294094338);
    Send_IMC_Command(32'd92570371);
    Send_IMC_Command(32'd293830660);
    Send_IMC_Command(32'd92372997);
    Send_IMC_Command(32'd293994502);
    Send_IMC_Command(32'd83952903);
    Send_IMC_Command(32'd293602056);
    Send_IMC_Command(32'd84018185);
    Send_IMC_Command(32'd84018442);
    Send_IMC_Command(32'd84083979);
    Send_IMC_Command(32'd293929740);
    Send_IMC_Command(32'd92700941);
    Send_IMC_Command(32'd293930766);
    Send_IMC_Command(32'd84151567);
    Send_IMC_Command(32'd92472848);
    Send_IMC_Command(32'd293962257);
    Send_IMC_Command(32'd293765394);
    Send_IMC_Command(32'd293962515);
    Send_IMC_Command(32'd92737812);
    Send_IMC_Command(32'd83955989);
    Send_IMC_Command(32'd84742934);
    Send_IMC_Command(32'd84087319);
    Send_IMC_Command(32'd84481816);
    Send_IMC_Command(32'd84480537);
    Send_IMC_Command(32'd84612634);
    Send_IMC_Command(32'd67769627);
    Send_IMC_Command(32'd67110428);
    Send_IMC_Command(32'd85531421);
    Send_IMC_Command(32'd67572766);
    Send_IMC_Command(32'd85859103);
    Send_IMC_Command(32'd67835424);
    Send_IMC_Command(32'd67176481);
    Send_IMC_Command(32'd85598242);
    Send_IMC_Command(32'd68095523);
    Send_IMC_Command(32'd86188068);
    Send_IMC_Command(32'd67311653);
    Send_IMC_Command(32'd68163366);
    Send_IMC_Command(32'd86385959);
    Send_IMC_Command(32'd67242280);
    Send_IMC_Command(32'd86517033);
    Send_IMC_Command(32'd85793834);
    Send_IMC_Command(32'd85918763);
    Send_IMC_Command(32'd86122796);
    Send_IMC_Command(32'd86255917);
    Send_IMC_Command(32'd86648622);
    Send_IMC_Command(32'd86714671);
    Send_IMC_Command(32'd86779696);
    Send_IMC_Command(32'd86838321);
    Send_IMC_Command(32'd87044402);
    Send_IMC_Command(32'd70266419);
    Send_IMC_Command(32'd86979380);
    Send_IMC_Command(32'd86912821);
    Send_IMC_Command(32'd87110454);
    Send_IMC_Command(32'd70661431);
    Send_IMC_Command(32'd70529592);
    Send_IMC_Command(32'd70136121);
    Send_IMC_Command(32'd70596922);
    Send_IMC_Command(32'd87372603);
    Send_IMC_Command(32'd70201404);
    Send_IMC_Command(32'd70401085);
    Send_IMC_Command(32'd87175998);
    Send_IMC_Command(32'd86980415);
    Send_IMC_Command(32'd87702336);
    Send_IMC_Command(32'd87111745);
    Send_IMC_Command(32'd87899714);
    Send_IMC_Command(32'd88097347);
    Send_IMC_Command(32'd88031556);
    Send_IMC_Command(32'd88031301);
    Send_IMC_Command(32'd88162886);
    Send_IMC_Command(32'd88359751);
    Send_IMC_Command(32'd71701832);
    Send_IMC_Command(32'd71435849);
    Send_IMC_Command(32'd71373898);
    Send_IMC_Command(32'd71636555);
    Send_IMC_Command(32'd71305292);
    Send_IMC_Command(32'd71241293);
    Send_IMC_Command(32'd71571534);
    Send_IMC_Command(32'd71767887);
    Send_IMC_Command(32'd71502160);
    Send_IMC_Command(32'd71699025);
    Send_IMC_Command(32'd71434322);
    Send_IMC_Command(32'd71370579);
    Send_IMC_Command(32'd71633748);
    Send_IMC_Command(32'd71303509);
    Send_IMC_Command(32'd71241558);
    Send_IMC_Command(32'd71566167);
    Send_IMC_Command(32'd71766104);
    Send_IMC_Command(32'd71500377);
    Send_IMC_Command(32'd89020250);
    Send_IMC_Command(32'd89412955);
    Send_IMC_Command(32'd89151580);
    Send_IMC_Command(32'd88689757);
    Send_IMC_Command(32'd88756830);
    Send_IMC_Command(32'd88624479);
    Send_IMC_Command(32'd88823392);
    Send_IMC_Command(32'd89807713);
    Send_IMC_Command(32'd88887138);
    Send_IMC_Command(32'd89217379);
    Send_IMC_Command(32'd89349732);
    Send_IMC_Command(32'd89808229);
    Send_IMC_Command(32'd88623718);
    Send_IMC_Command(32'd88821095);
    Send_IMC_Command(32'd88823912);
    Send_IMC_Command(32'd89150825);
    Send_IMC_Command(32'd89347946);
    Send_IMC_Command(32'd89414763);
    Send_IMC_Command(32'd89743212);
    Send_IMC_Command(32'd89939309);
    Send_IMC_Command(32'd90071150);
    Send_IMC_Command(32'd89940335);
    Send_IMC_Command(32'd90268272);
    Send_IMC_Command(32'd90136945);
    Send_IMC_Command(32'd90203250);
    Send_IMC_Command(32'd90400115);
    Send_IMC_Command(32'd90467444);
    Send_IMC_Command(32'd90534517);
    Send_IMC_Command(32'd90795638);
    Send_IMC_Command(32'd90664839);
    Send_IMC_Command(32'd91453062);
    Send_IMC_Command(32'd90928517);
    Send_IMC_Command(32'd90599300);
    Send_IMC_Command(32'd91255939);
    Send_IMC_Command(32'd91058562);
    Send_IMC_Command(32'd90730625);
    Send_IMC_Command(32'd90401408);
    Send_IMC_Command(32'd93293568);
    Send_IMC_Command(32'd294554625);
    Send_IMC_Command(32'd294620674);
    Send_IMC_Command(32'd93096707);
    Send_IMC_Command(32'd294356996);
    Send_IMC_Command(32'd92899333);
    Send_IMC_Command(32'd294518790);
    Send_IMC_Command(32'd83952903);
    Send_IMC_Command(32'd294126344);
    Send_IMC_Command(32'd84018185);
    Send_IMC_Command(32'd84018442);
    Send_IMC_Command(32'd84083979);
    Send_IMC_Command(32'd294454028);
    Send_IMC_Command(32'd93227277);
    Send_IMC_Command(32'd294455054);
    Send_IMC_Command(32'd84151567);
    Send_IMC_Command(32'd92997136);
    Send_IMC_Command(32'd294488593);
    Send_IMC_Command(32'd294291730);
    Send_IMC_Command(32'd294488851);
    Send_IMC_Command(32'd93262100);
    Send_IMC_Command(32'd83955989);
    Send_IMC_Command(32'd84742934);
    Send_IMC_Command(32'd84087319);
    Send_IMC_Command(32'd84481816);
    Send_IMC_Command(32'd84480537);
    Send_IMC_Command(32'd84612634);
    Send_IMC_Command(32'd67769627);
    Send_IMC_Command(32'd67110428);
    Send_IMC_Command(32'd85531421);
    Send_IMC_Command(32'd67572766);
    Send_IMC_Command(32'd85859103);
    Send_IMC_Command(32'd67835424);
    Send_IMC_Command(32'd67176481);
    Send_IMC_Command(32'd85598242);
    Send_IMC_Command(32'd68095523);
    Send_IMC_Command(32'd86188068);
    Send_IMC_Command(32'd67311653);
    Send_IMC_Command(32'd68163366);
    Send_IMC_Command(32'd86385959);
    Send_IMC_Command(32'd67242280);
    Send_IMC_Command(32'd86517033);
    Send_IMC_Command(32'd85793834);
    Send_IMC_Command(32'd85918763);
    Send_IMC_Command(32'd86122796);
    Send_IMC_Command(32'd86255917);
    Send_IMC_Command(32'd86648622);
    Send_IMC_Command(32'd86714671);
    Send_IMC_Command(32'd86779696);
    Send_IMC_Command(32'd86838321);
    Send_IMC_Command(32'd87044402);
    Send_IMC_Command(32'd70266419);
    Send_IMC_Command(32'd86979380);
    Send_IMC_Command(32'd86912821);
    Send_IMC_Command(32'd87110454);
    Send_IMC_Command(32'd70661431);
    Send_IMC_Command(32'd70529592);
    Send_IMC_Command(32'd70136121);
    Send_IMC_Command(32'd70596922);
    Send_IMC_Command(32'd87372603);
    Send_IMC_Command(32'd70201404);
    Send_IMC_Command(32'd70401085);
    Send_IMC_Command(32'd87175998);
    Send_IMC_Command(32'd86980415);
    Send_IMC_Command(32'd87702336);
    Send_IMC_Command(32'd87111745);
    Send_IMC_Command(32'd87899714);
    Send_IMC_Command(32'd88097347);
    Send_IMC_Command(32'd88031556);
    Send_IMC_Command(32'd88031301);
    Send_IMC_Command(32'd88162886);
    Send_IMC_Command(32'd88359751);
    Send_IMC_Command(32'd71701832);
    Send_IMC_Command(32'd71435849);
    Send_IMC_Command(32'd71373898);
    Send_IMC_Command(32'd71636555);
    Send_IMC_Command(32'd71305292);
    Send_IMC_Command(32'd71241293);
    Send_IMC_Command(32'd71571534);
    Send_IMC_Command(32'd71767887);
    Send_IMC_Command(32'd71502160);
    Send_IMC_Command(32'd71699025);
    Send_IMC_Command(32'd71434322);
    Send_IMC_Command(32'd71370579);
    Send_IMC_Command(32'd71633748);
    Send_IMC_Command(32'd71303509);
    Send_IMC_Command(32'd71241558);
    Send_IMC_Command(32'd71566167);
    Send_IMC_Command(32'd71766104);
    Send_IMC_Command(32'd71500377);
    Send_IMC_Command(32'd89020250);
    Send_IMC_Command(32'd89412955);
    Send_IMC_Command(32'd89151580);
    Send_IMC_Command(32'd88689757);
    Send_IMC_Command(32'd88756830);
    Send_IMC_Command(32'd88624479);
    Send_IMC_Command(32'd88823392);
    Send_IMC_Command(32'd89807713);
    Send_IMC_Command(32'd88887138);
    Send_IMC_Command(32'd89217379);
    Send_IMC_Command(32'd89349732);
    Send_IMC_Command(32'd89808229);
    Send_IMC_Command(32'd88623718);
    Send_IMC_Command(32'd88821095);
    Send_IMC_Command(32'd88823912);
    Send_IMC_Command(32'd89150825);
    Send_IMC_Command(32'd89347946);
    Send_IMC_Command(32'd89414763);
    Send_IMC_Command(32'd89743212);
    Send_IMC_Command(32'd89939309);
    Send_IMC_Command(32'd90071150);
    Send_IMC_Command(32'd89940335);
    Send_IMC_Command(32'd90268272);
    Send_IMC_Command(32'd90136945);
    Send_IMC_Command(32'd90203250);
    Send_IMC_Command(32'd90400115);
    Send_IMC_Command(32'd90467444);
    Send_IMC_Command(32'd90534517);
    Send_IMC_Command(32'd90795638);
    Send_IMC_Command(32'd90664847);
    Send_IMC_Command(32'd91453070);
    Send_IMC_Command(32'd90928525);
    Send_IMC_Command(32'd90599308);
    Send_IMC_Command(32'd91255947);
    Send_IMC_Command(32'd91058570);
    Send_IMC_Command(32'd90730633);
    Send_IMC_Command(32'd90401416);
    Send_IMC_Command(32'd93819904);
    Send_IMC_Command(32'd295080961);
    Send_IMC_Command(32'd295147010);
    Send_IMC_Command(32'd93623043);
    Send_IMC_Command(32'd294883332);
    Send_IMC_Command(32'd93425669);
    Send_IMC_Command(32'd295043078);
    Send_IMC_Command(32'd83952903);
    Send_IMC_Command(32'd294650632);
    Send_IMC_Command(32'd84018185);
    Send_IMC_Command(32'd84018442);
    Send_IMC_Command(32'd84083979);
    Send_IMC_Command(32'd294978316);
    Send_IMC_Command(32'd93753613);
    Send_IMC_Command(32'd294979342);
    Send_IMC_Command(32'd84151567);
    Send_IMC_Command(32'd93521424);
    Send_IMC_Command(32'd295014929);
    Send_IMC_Command(32'd294818066);
    Send_IMC_Command(32'd295015187);
    Send_IMC_Command(32'd93786388);
    Send_IMC_Command(32'd83955989);
    Send_IMC_Command(32'd84742934);
    Send_IMC_Command(32'd84087319);
    Send_IMC_Command(32'd84481816);
    Send_IMC_Command(32'd84480537);
    Send_IMC_Command(32'd84612634);
    Send_IMC_Command(32'd67769627);
    Send_IMC_Command(32'd67110428);
    Send_IMC_Command(32'd85531421);
    Send_IMC_Command(32'd67572766);
    Send_IMC_Command(32'd85859103);
    Send_IMC_Command(32'd67835424);
    Send_IMC_Command(32'd67176481);
    Send_IMC_Command(32'd85598242);
    Send_IMC_Command(32'd68095523);
    Send_IMC_Command(32'd86188068);
    Send_IMC_Command(32'd67311653);
    Send_IMC_Command(32'd68163366);
    Send_IMC_Command(32'd86385959);
    Send_IMC_Command(32'd67242280);
    Send_IMC_Command(32'd86517033);
    Send_IMC_Command(32'd85793834);
    Send_IMC_Command(32'd85918763);
    Send_IMC_Command(32'd86122796);
    Send_IMC_Command(32'd86255917);
    Send_IMC_Command(32'd86648622);
    Send_IMC_Command(32'd86714671);
    Send_IMC_Command(32'd86779696);
    Send_IMC_Command(32'd86838321);
    Send_IMC_Command(32'd87044402);
    Send_IMC_Command(32'd70266419);
    Send_IMC_Command(32'd86979380);
    Send_IMC_Command(32'd86912821);
    Send_IMC_Command(32'd87110454);
    Send_IMC_Command(32'd70661431);
    Send_IMC_Command(32'd70529592);
    Send_IMC_Command(32'd70136121);
    Send_IMC_Command(32'd70596922);
    Send_IMC_Command(32'd87372603);
    Send_IMC_Command(32'd70201404);
    Send_IMC_Command(32'd70401085);
    Send_IMC_Command(32'd87175998);
    Send_IMC_Command(32'd86980415);
    Send_IMC_Command(32'd87702336);
    Send_IMC_Command(32'd87111745);
    Send_IMC_Command(32'd87899714);
    Send_IMC_Command(32'd88097347);
    Send_IMC_Command(32'd88031556);
    Send_IMC_Command(32'd88031301);
    Send_IMC_Command(32'd88162886);
    Send_IMC_Command(32'd88359751);
    Send_IMC_Command(32'd71701832);
    Send_IMC_Command(32'd71435849);
    Send_IMC_Command(32'd71373898);
    Send_IMC_Command(32'd71636555);
    Send_IMC_Command(32'd71305292);
    Send_IMC_Command(32'd71241293);
    Send_IMC_Command(32'd71571534);
    Send_IMC_Command(32'd71767887);
    Send_IMC_Command(32'd71502160);
    Send_IMC_Command(32'd71699025);
    Send_IMC_Command(32'd71434322);
    Send_IMC_Command(32'd71370579);
    Send_IMC_Command(32'd71633748);
    Send_IMC_Command(32'd71303509);
    Send_IMC_Command(32'd71241558);
    Send_IMC_Command(32'd71566167);
    Send_IMC_Command(32'd71766104);
    Send_IMC_Command(32'd71500377);
    Send_IMC_Command(32'd89020250);
    Send_IMC_Command(32'd89412955);
    Send_IMC_Command(32'd89151580);
    Send_IMC_Command(32'd88689757);
    Send_IMC_Command(32'd88756830);
    Send_IMC_Command(32'd88624479);
    Send_IMC_Command(32'd88823392);
    Send_IMC_Command(32'd89807713);
    Send_IMC_Command(32'd88887138);
    Send_IMC_Command(32'd89217379);
    Send_IMC_Command(32'd89349732);
    Send_IMC_Command(32'd89808229);
    Send_IMC_Command(32'd88623718);
    Send_IMC_Command(32'd88821095);
    Send_IMC_Command(32'd88823912);
    Send_IMC_Command(32'd89150825);
    Send_IMC_Command(32'd89347946);
    Send_IMC_Command(32'd89414763);
    Send_IMC_Command(32'd89743212);
    Send_IMC_Command(32'd89939309);
    Send_IMC_Command(32'd90071150);
    Send_IMC_Command(32'd89940335);
    Send_IMC_Command(32'd90268272);
    Send_IMC_Command(32'd90136945);
    Send_IMC_Command(32'd90203250);
    Send_IMC_Command(32'd90400115);
    Send_IMC_Command(32'd90467444);
    Send_IMC_Command(32'd90534517);
    Send_IMC_Command(32'd90795638);
    Send_IMC_Command(32'd90664855);
    Send_IMC_Command(32'd91453078);
    Send_IMC_Command(32'd90928533);
    Send_IMC_Command(32'd90599316);
    Send_IMC_Command(32'd91255955);
    Send_IMC_Command(32'd91058578);
    Send_IMC_Command(32'd90730641);
    Send_IMC_Command(32'd90401424);
    Send_IMC_Command(32'd94346240);
    Send_IMC_Command(32'd295607297);
    Send_IMC_Command(32'd295673346);
    Send_IMC_Command(32'd94149379);
    Send_IMC_Command(32'd295409668);
    Send_IMC_Command(32'd93952005);
    Send_IMC_Command(32'd295567366);
    Send_IMC_Command(32'd83952903);
    Send_IMC_Command(32'd295174920);
    Send_IMC_Command(32'd84018185);
    Send_IMC_Command(32'd84018442);
    Send_IMC_Command(32'd84083979);
    Send_IMC_Command(32'd295502604);
    Send_IMC_Command(32'd94279949);
    Send_IMC_Command(32'd295503630);
    Send_IMC_Command(32'd84151567);
    Send_IMC_Command(32'd94045712);
    Send_IMC_Command(32'd295541265);
    Send_IMC_Command(32'd295344402);
    Send_IMC_Command(32'd295541523);
    Send_IMC_Command(32'd94310676);
    Send_IMC_Command(32'd83955989);
    Send_IMC_Command(32'd84742934);
    Send_IMC_Command(32'd84087319);
    Send_IMC_Command(32'd84481816);
    Send_IMC_Command(32'd84480537);
    Send_IMC_Command(32'd84612634);
    Send_IMC_Command(32'd67769627);
    Send_IMC_Command(32'd67110428);
    Send_IMC_Command(32'd85531421);
    Send_IMC_Command(32'd67572766);
    Send_IMC_Command(32'd85859103);
    Send_IMC_Command(32'd67835424);
    Send_IMC_Command(32'd67176481);
    Send_IMC_Command(32'd85598242);
    Send_IMC_Command(32'd68095523);
    Send_IMC_Command(32'd86188068);
    Send_IMC_Command(32'd67311653);
    Send_IMC_Command(32'd68163366);
    Send_IMC_Command(32'd86385959);
    Send_IMC_Command(32'd67242280);
    Send_IMC_Command(32'd86517033);
    Send_IMC_Command(32'd85793834);
    Send_IMC_Command(32'd85918763);
    Send_IMC_Command(32'd86122796);
    Send_IMC_Command(32'd86255917);
    Send_IMC_Command(32'd86648622);
    Send_IMC_Command(32'd86714671);
    Send_IMC_Command(32'd86779696);
    Send_IMC_Command(32'd86838321);
    Send_IMC_Command(32'd87044402);
    Send_IMC_Command(32'd70266419);
    Send_IMC_Command(32'd86979380);
    Send_IMC_Command(32'd86912821);
    Send_IMC_Command(32'd87110454);
    Send_IMC_Command(32'd70661431);
    Send_IMC_Command(32'd70529592);
    Send_IMC_Command(32'd70136121);
    Send_IMC_Command(32'd70596922);
    Send_IMC_Command(32'd87372603);
    Send_IMC_Command(32'd70201404);
    Send_IMC_Command(32'd70401085);
    Send_IMC_Command(32'd87175998);
    Send_IMC_Command(32'd86980415);
    Send_IMC_Command(32'd87702336);
    Send_IMC_Command(32'd87111745);
    Send_IMC_Command(32'd87899714);
    Send_IMC_Command(32'd88097347);
    Send_IMC_Command(32'd88031556);
    Send_IMC_Command(32'd88031301);
    Send_IMC_Command(32'd88162886);
    Send_IMC_Command(32'd88359751);
    Send_IMC_Command(32'd71701832);
    Send_IMC_Command(32'd71435849);
    Send_IMC_Command(32'd71373898);
    Send_IMC_Command(32'd71636555);
    Send_IMC_Command(32'd71305292);
    Send_IMC_Command(32'd71241293);
    Send_IMC_Command(32'd71571534);
    Send_IMC_Command(32'd71767887);
    Send_IMC_Command(32'd71502160);
    Send_IMC_Command(32'd71699025);
    Send_IMC_Command(32'd71434322);
    Send_IMC_Command(32'd71370579);
    Send_IMC_Command(32'd71633748);
    Send_IMC_Command(32'd71303509);
    Send_IMC_Command(32'd71241558);
    Send_IMC_Command(32'd71566167);
    Send_IMC_Command(32'd71766104);
    Send_IMC_Command(32'd71500377);
    Send_IMC_Command(32'd89020250);
    Send_IMC_Command(32'd89412955);
    Send_IMC_Command(32'd89151580);
    Send_IMC_Command(32'd88689757);
    Send_IMC_Command(32'd88756830);
    Send_IMC_Command(32'd88624479);
    Send_IMC_Command(32'd88823392);
    Send_IMC_Command(32'd89807713);
    Send_IMC_Command(32'd88887138);
    Send_IMC_Command(32'd89217379);
    Send_IMC_Command(32'd89349732);
    Send_IMC_Command(32'd89808229);
    Send_IMC_Command(32'd88623718);
    Send_IMC_Command(32'd88821095);
    Send_IMC_Command(32'd88823912);
    Send_IMC_Command(32'd89150825);
    Send_IMC_Command(32'd89347946);
    Send_IMC_Command(32'd89414763);
    Send_IMC_Command(32'd89743212);
    Send_IMC_Command(32'd89939309);
    Send_IMC_Command(32'd90071150);
    Send_IMC_Command(32'd89940335);
    Send_IMC_Command(32'd90268272);
    Send_IMC_Command(32'd90136945);
    Send_IMC_Command(32'd90203250);
    Send_IMC_Command(32'd90400115);
    Send_IMC_Command(32'd90467444);
    Send_IMC_Command(32'd90534517);
    Send_IMC_Command(32'd90795638);
    Send_IMC_Command(32'd90664863);
    Send_IMC_Command(32'd91453086);
    Send_IMC_Command(32'd90928541);
    Send_IMC_Command(32'd90599324);
    Send_IMC_Command(32'd91255963);
    Send_IMC_Command(32'd91058586);
    Send_IMC_Command(32'd90730649);
    Send_IMC_Command(32'd90401432);
    Send_IMC_Command(32'd94872576);
    Send_IMC_Command(32'd296133633);
    Send_IMC_Command(32'd296199682);
    Send_IMC_Command(32'd94675715);
    Send_IMC_Command(32'd295936004);
    Send_IMC_Command(32'd94478341);
    Send_IMC_Command(32'd296091654);
    Send_IMC_Command(32'd83952903);
    Send_IMC_Command(32'd295699208);
    Send_IMC_Command(32'd84018185);
    Send_IMC_Command(32'd84018442);
    Send_IMC_Command(32'd84083979);
    Send_IMC_Command(32'd296026892);
    Send_IMC_Command(32'd94806285);
    Send_IMC_Command(32'd296027918);
    Send_IMC_Command(32'd84151567);
    Send_IMC_Command(32'd94570000);
    Send_IMC_Command(32'd296067601);
    Send_IMC_Command(32'd295870738);
    Send_IMC_Command(32'd296067859);
    Send_IMC_Command(32'd94834964);
    Send_IMC_Command(32'd83955989);
    Send_IMC_Command(32'd84742934);
    Send_IMC_Command(32'd84087319);
    Send_IMC_Command(32'd84481816);
    Send_IMC_Command(32'd84480537);
    Send_IMC_Command(32'd84612634);
    Send_IMC_Command(32'd67769627);
    Send_IMC_Command(32'd67110428);
    Send_IMC_Command(32'd85531421);
    Send_IMC_Command(32'd67572766);
    Send_IMC_Command(32'd85859103);
    Send_IMC_Command(32'd67835424);
    Send_IMC_Command(32'd67176481);
    Send_IMC_Command(32'd85598242);
    Send_IMC_Command(32'd68095523);
    Send_IMC_Command(32'd86188068);
    Send_IMC_Command(32'd67311653);
    Send_IMC_Command(32'd68163366);
    Send_IMC_Command(32'd86385959);
    Send_IMC_Command(32'd67242280);
    Send_IMC_Command(32'd86517033);
    Send_IMC_Command(32'd85793834);
    Send_IMC_Command(32'd85918763);
    Send_IMC_Command(32'd86122796);
    Send_IMC_Command(32'd86255917);
    Send_IMC_Command(32'd86648622);
    Send_IMC_Command(32'd86714671);
    Send_IMC_Command(32'd86779696);
    Send_IMC_Command(32'd86838321);
    Send_IMC_Command(32'd87044402);
    Send_IMC_Command(32'd70266419);
    Send_IMC_Command(32'd86979380);
    Send_IMC_Command(32'd86912821);
    Send_IMC_Command(32'd87110454);
    Send_IMC_Command(32'd70661431);
    Send_IMC_Command(32'd70529592);
    Send_IMC_Command(32'd70136121);
    Send_IMC_Command(32'd70596922);
    Send_IMC_Command(32'd87372603);
    Send_IMC_Command(32'd70201404);
    Send_IMC_Command(32'd70401085);
    Send_IMC_Command(32'd87175998);
    Send_IMC_Command(32'd86980415);
    Send_IMC_Command(32'd87702336);
    Send_IMC_Command(32'd87111745);
    Send_IMC_Command(32'd87899714);
    Send_IMC_Command(32'd88097347);
    Send_IMC_Command(32'd88031556);
    Send_IMC_Command(32'd88031301);
    Send_IMC_Command(32'd88162886);
    Send_IMC_Command(32'd88359751);
    Send_IMC_Command(32'd71701832);
    Send_IMC_Command(32'd71435849);
    Send_IMC_Command(32'd71373898);
    Send_IMC_Command(32'd71636555);
    Send_IMC_Command(32'd71305292);
    Send_IMC_Command(32'd71241293);
    Send_IMC_Command(32'd71571534);
    Send_IMC_Command(32'd71767887);
    Send_IMC_Command(32'd71502160);
    Send_IMC_Command(32'd71699025);
    Send_IMC_Command(32'd71434322);
    Send_IMC_Command(32'd71370579);
    Send_IMC_Command(32'd71633748);
    Send_IMC_Command(32'd71303509);
    Send_IMC_Command(32'd71241558);
    Send_IMC_Command(32'd71566167);
    Send_IMC_Command(32'd71766104);
    Send_IMC_Command(32'd71500377);
    Send_IMC_Command(32'd89020250);
    Send_IMC_Command(32'd89412955);
    Send_IMC_Command(32'd89151580);
    Send_IMC_Command(32'd88689757);
    Send_IMC_Command(32'd88756830);
    Send_IMC_Command(32'd88624479);
    Send_IMC_Command(32'd88823392);
    Send_IMC_Command(32'd89807713);
    Send_IMC_Command(32'd88887138);
    Send_IMC_Command(32'd89217379);
    Send_IMC_Command(32'd89349732);
    Send_IMC_Command(32'd89808229);
    Send_IMC_Command(32'd88623718);
    Send_IMC_Command(32'd88821095);
    Send_IMC_Command(32'd88823912);
    Send_IMC_Command(32'd89150825);
    Send_IMC_Command(32'd89347946);
    Send_IMC_Command(32'd89414763);
    Send_IMC_Command(32'd89743212);
    Send_IMC_Command(32'd89939309);
    Send_IMC_Command(32'd90071150);
    Send_IMC_Command(32'd89940335);
    Send_IMC_Command(32'd90268272);
    Send_IMC_Command(32'd90136945);
    Send_IMC_Command(32'd90203250);
    Send_IMC_Command(32'd90400115);
    Send_IMC_Command(32'd90467444);
    Send_IMC_Command(32'd90534517);
    Send_IMC_Command(32'd90795638);
    Send_IMC_Command(32'd90664871);
    Send_IMC_Command(32'd91453094);
    Send_IMC_Command(32'd90928549);
    Send_IMC_Command(32'd90599332);
    Send_IMC_Command(32'd91255971);
    Send_IMC_Command(32'd91058594);
    Send_IMC_Command(32'd90730657);
    Send_IMC_Command(32'd90401440);
    Send_IMC_Command(32'd95398912);
    Send_IMC_Command(32'd296659969);
    Send_IMC_Command(32'd296726018);
    Send_IMC_Command(32'd95202051);
    Send_IMC_Command(32'd296462340);
    Send_IMC_Command(32'd95004677);
    Send_IMC_Command(32'd296615942);
    Send_IMC_Command(32'd83952903);
    Send_IMC_Command(32'd296223496);
    Send_IMC_Command(32'd84018185);
    Send_IMC_Command(32'd84018442);
    Send_IMC_Command(32'd84083979);
    Send_IMC_Command(32'd296551180);
    Send_IMC_Command(32'd95332621);
    Send_IMC_Command(32'd296552206);
    Send_IMC_Command(32'd84151567);
    Send_IMC_Command(32'd95094288);
    Send_IMC_Command(32'd296593937);
    Send_IMC_Command(32'd296397074);
    Send_IMC_Command(32'd296594195);
    Send_IMC_Command(32'd95359252);
    Send_IMC_Command(32'd83955989);
    Send_IMC_Command(32'd84742934);
    Send_IMC_Command(32'd84087319);
    Send_IMC_Command(32'd84481816);
    Send_IMC_Command(32'd84480537);
    Send_IMC_Command(32'd84612634);
    Send_IMC_Command(32'd67769627);
    Send_IMC_Command(32'd67110428);
    Send_IMC_Command(32'd85531421);
    Send_IMC_Command(32'd67572766);
    Send_IMC_Command(32'd85859103);
    Send_IMC_Command(32'd67835424);
    Send_IMC_Command(32'd67176481);
    Send_IMC_Command(32'd85598242);
    Send_IMC_Command(32'd68095523);
    Send_IMC_Command(32'd86188068);
    Send_IMC_Command(32'd67311653);
    Send_IMC_Command(32'd68163366);
    Send_IMC_Command(32'd86385959);
    Send_IMC_Command(32'd67242280);
    Send_IMC_Command(32'd86517033);
    Send_IMC_Command(32'd85793834);
    Send_IMC_Command(32'd85918763);
    Send_IMC_Command(32'd86122796);
    Send_IMC_Command(32'd86255917);
    Send_IMC_Command(32'd86648622);
    Send_IMC_Command(32'd86714671);
    Send_IMC_Command(32'd86779696);
    Send_IMC_Command(32'd86838321);
    Send_IMC_Command(32'd87044402);
    Send_IMC_Command(32'd70266419);
    Send_IMC_Command(32'd86979380);
    Send_IMC_Command(32'd86912821);
    Send_IMC_Command(32'd87110454);
    Send_IMC_Command(32'd70661431);
    Send_IMC_Command(32'd70529592);
    Send_IMC_Command(32'd70136121);
    Send_IMC_Command(32'd70596922);
    Send_IMC_Command(32'd87372603);
    Send_IMC_Command(32'd70201404);
    Send_IMC_Command(32'd70401085);
    Send_IMC_Command(32'd87175998);
    Send_IMC_Command(32'd86980415);
    Send_IMC_Command(32'd87702336);
    Send_IMC_Command(32'd87111745);
    Send_IMC_Command(32'd87899714);
    Send_IMC_Command(32'd88097347);
    Send_IMC_Command(32'd88031556);
    Send_IMC_Command(32'd88031301);
    Send_IMC_Command(32'd88162886);
    Send_IMC_Command(32'd88359751);
    Send_IMC_Command(32'd71701832);
    Send_IMC_Command(32'd71435849);
    Send_IMC_Command(32'd71373898);
    Send_IMC_Command(32'd71636555);
    Send_IMC_Command(32'd71305292);
    Send_IMC_Command(32'd71241293);
    Send_IMC_Command(32'd71571534);
    Send_IMC_Command(32'd71767887);
    Send_IMC_Command(32'd71502160);
    Send_IMC_Command(32'd71699025);
    Send_IMC_Command(32'd71434322);
    Send_IMC_Command(32'd71370579);
    Send_IMC_Command(32'd71633748);
    Send_IMC_Command(32'd71303509);
    Send_IMC_Command(32'd71241558);
    Send_IMC_Command(32'd71566167);
    Send_IMC_Command(32'd71766104);
    Send_IMC_Command(32'd71500377);
    Send_IMC_Command(32'd89020250);
    Send_IMC_Command(32'd89412955);
    Send_IMC_Command(32'd89151580);
    Send_IMC_Command(32'd88689757);
    Send_IMC_Command(32'd88756830);
    Send_IMC_Command(32'd88624479);
    Send_IMC_Command(32'd88823392);
    Send_IMC_Command(32'd89807713);
    Send_IMC_Command(32'd88887138);
    Send_IMC_Command(32'd89217379);
    Send_IMC_Command(32'd89349732);
    Send_IMC_Command(32'd89808229);
    Send_IMC_Command(32'd88623718);
    Send_IMC_Command(32'd88821095);
    Send_IMC_Command(32'd88823912);
    Send_IMC_Command(32'd89150825);
    Send_IMC_Command(32'd89347946);
    Send_IMC_Command(32'd89414763);
    Send_IMC_Command(32'd89743212);
    Send_IMC_Command(32'd89939309);
    Send_IMC_Command(32'd90071150);
    Send_IMC_Command(32'd89940335);
    Send_IMC_Command(32'd90268272);
    Send_IMC_Command(32'd90136945);
    Send_IMC_Command(32'd90203250);
    Send_IMC_Command(32'd90400115);
    Send_IMC_Command(32'd90467444);
    Send_IMC_Command(32'd90534517);
    Send_IMC_Command(32'd90795638);
    Send_IMC_Command(32'd90664879);
    Send_IMC_Command(32'd91453102);
    Send_IMC_Command(32'd90928557);
    Send_IMC_Command(32'd90599340);
    Send_IMC_Command(32'd91255979);
    Send_IMC_Command(32'd91058602);
    Send_IMC_Command(32'd90730665);
    Send_IMC_Command(32'd90401448);
    Send_IMC_Command(32'd95925248);
    Send_IMC_Command(32'd297186305);
    Send_IMC_Command(32'd297252354);
    Send_IMC_Command(32'd95728387);
    Send_IMC_Command(32'd296988676);
    Send_IMC_Command(32'd95531013);
    Send_IMC_Command(32'd297140230);
    Send_IMC_Command(32'd83952903);
    Send_IMC_Command(32'd296747784);
    Send_IMC_Command(32'd84018185);
    Send_IMC_Command(32'd84018442);
    Send_IMC_Command(32'd84083979);
    Send_IMC_Command(32'd297075468);
    Send_IMC_Command(32'd95858957);
    Send_IMC_Command(32'd297076494);
    Send_IMC_Command(32'd84151567);
    Send_IMC_Command(32'd95618576);
    Send_IMC_Command(32'd297120273);
    Send_IMC_Command(32'd296923410);
    Send_IMC_Command(32'd297120531);
    Send_IMC_Command(32'd95883540);
    Send_IMC_Command(32'd83955989);
    Send_IMC_Command(32'd84742934);
    Send_IMC_Command(32'd84087319);
    Send_IMC_Command(32'd84481816);
    Send_IMC_Command(32'd84480537);
    Send_IMC_Command(32'd84612634);
    Send_IMC_Command(32'd67769627);
    Send_IMC_Command(32'd67110428);
    Send_IMC_Command(32'd85531421);
    Send_IMC_Command(32'd67572766);
    Send_IMC_Command(32'd85859103);
    Send_IMC_Command(32'd67835424);
    Send_IMC_Command(32'd67176481);
    Send_IMC_Command(32'd85598242);
    Send_IMC_Command(32'd68095523);
    Send_IMC_Command(32'd86188068);
    Send_IMC_Command(32'd67311653);
    Send_IMC_Command(32'd68163366);
    Send_IMC_Command(32'd86385959);
    Send_IMC_Command(32'd67242280);
    Send_IMC_Command(32'd86517033);
    Send_IMC_Command(32'd85793834);
    Send_IMC_Command(32'd85918763);
    Send_IMC_Command(32'd86122796);
    Send_IMC_Command(32'd86255917);
    Send_IMC_Command(32'd86648622);
    Send_IMC_Command(32'd86714671);
    Send_IMC_Command(32'd86779696);
    Send_IMC_Command(32'd86838321);
    Send_IMC_Command(32'd87044402);
    Send_IMC_Command(32'd70266419);
    Send_IMC_Command(32'd86979380);
    Send_IMC_Command(32'd86912821);
    Send_IMC_Command(32'd87110454);
    Send_IMC_Command(32'd70661431);
    Send_IMC_Command(32'd70529592);
    Send_IMC_Command(32'd70136121);
    Send_IMC_Command(32'd70596922);
    Send_IMC_Command(32'd87372603);
    Send_IMC_Command(32'd70201404);
    Send_IMC_Command(32'd70401085);
    Send_IMC_Command(32'd87175998);
    Send_IMC_Command(32'd86980415);
    Send_IMC_Command(32'd87702336);
    Send_IMC_Command(32'd87111745);
    Send_IMC_Command(32'd87899714);
    Send_IMC_Command(32'd88097347);
    Send_IMC_Command(32'd88031556);
    Send_IMC_Command(32'd88031301);
    Send_IMC_Command(32'd88162886);
    Send_IMC_Command(32'd88359751);
    Send_IMC_Command(32'd71701832);
    Send_IMC_Command(32'd71435849);
    Send_IMC_Command(32'd71373898);
    Send_IMC_Command(32'd71636555);
    Send_IMC_Command(32'd71305292);
    Send_IMC_Command(32'd71241293);
    Send_IMC_Command(32'd71571534);
    Send_IMC_Command(32'd71767887);
    Send_IMC_Command(32'd71502160);
    Send_IMC_Command(32'd71699025);
    Send_IMC_Command(32'd71434322);
    Send_IMC_Command(32'd71370579);
    Send_IMC_Command(32'd71633748);
    Send_IMC_Command(32'd71303509);
    Send_IMC_Command(32'd71241558);
    Send_IMC_Command(32'd71566167);
    Send_IMC_Command(32'd71766104);
    Send_IMC_Command(32'd71500377);
    Send_IMC_Command(32'd89020250);
    Send_IMC_Command(32'd89412955);
    Send_IMC_Command(32'd89151580);
    Send_IMC_Command(32'd88689757);
    Send_IMC_Command(32'd88756830);
    Send_IMC_Command(32'd88624479);
    Send_IMC_Command(32'd88823392);
    Send_IMC_Command(32'd89807713);
    Send_IMC_Command(32'd88887138);
    Send_IMC_Command(32'd89217379);
    Send_IMC_Command(32'd89349732);
    Send_IMC_Command(32'd89808229);
    Send_IMC_Command(32'd88623718);
    Send_IMC_Command(32'd88821095);
    Send_IMC_Command(32'd88823912);
    Send_IMC_Command(32'd89150825);
    Send_IMC_Command(32'd89347946);
    Send_IMC_Command(32'd89414763);
    Send_IMC_Command(32'd89743212);
    Send_IMC_Command(32'd89939309);
    Send_IMC_Command(32'd90071150);
    Send_IMC_Command(32'd89940335);
    Send_IMC_Command(32'd90268272);
    Send_IMC_Command(32'd90136945);
    Send_IMC_Command(32'd90203250);
    Send_IMC_Command(32'd90400115);
    Send_IMC_Command(32'd90467444);
    Send_IMC_Command(32'd90534517);
    Send_IMC_Command(32'd90795638);
    Send_IMC_Command(32'd90664887);
    Send_IMC_Command(32'd91453110);
    Send_IMC_Command(32'd90928565);
    Send_IMC_Command(32'd90599348);
    Send_IMC_Command(32'd91255987);
    Send_IMC_Command(32'd91058610);
    Send_IMC_Command(32'd90730673);
    Send_IMC_Command(32'd90401456);
    Send_IMC_Command(32'd96451584);
    Send_IMC_Command(32'd297712641);
    Send_IMC_Command(32'd297778690);
    Send_IMC_Command(32'd96254723);
    Send_IMC_Command(32'd297515012);
    Send_IMC_Command(32'd96057349);
    Send_IMC_Command(32'd297664518);
    Send_IMC_Command(32'd83952903);
    Send_IMC_Command(32'd297272072);
    Send_IMC_Command(32'd84018185);
    Send_IMC_Command(32'd84018442);
    Send_IMC_Command(32'd84083979);
    Send_IMC_Command(32'd297599756);
    Send_IMC_Command(32'd96385293);
    Send_IMC_Command(32'd297600782);
    Send_IMC_Command(32'd84151567);
    Send_IMC_Command(32'd96142864);
    Send_IMC_Command(32'd297646609);
    Send_IMC_Command(32'd297449746);
    Send_IMC_Command(32'd297646867);
    Send_IMC_Command(32'd96407828);
    Send_IMC_Command(32'd83955989);
    Send_IMC_Command(32'd84742934);
    Send_IMC_Command(32'd84087319);
    Send_IMC_Command(32'd84481816);
    Send_IMC_Command(32'd84480537);
    Send_IMC_Command(32'd84612634);
    Send_IMC_Command(32'd67769627);
    Send_IMC_Command(32'd67110428);
    Send_IMC_Command(32'd85531421);
    Send_IMC_Command(32'd67572766);
    Send_IMC_Command(32'd85859103);
    Send_IMC_Command(32'd67835424);
    Send_IMC_Command(32'd67176481);
    Send_IMC_Command(32'd85598242);
    Send_IMC_Command(32'd68095523);
    Send_IMC_Command(32'd86188068);
    Send_IMC_Command(32'd67311653);
    Send_IMC_Command(32'd68163366);
    Send_IMC_Command(32'd86385959);
    Send_IMC_Command(32'd67242280);
    Send_IMC_Command(32'd86517033);
    Send_IMC_Command(32'd85793834);
    Send_IMC_Command(32'd85918763);
    Send_IMC_Command(32'd86122796);
    Send_IMC_Command(32'd86255917);
    Send_IMC_Command(32'd86648622);
    Send_IMC_Command(32'd86714671);
    Send_IMC_Command(32'd86779696);
    Send_IMC_Command(32'd86838321);
    Send_IMC_Command(32'd87044402);
    Send_IMC_Command(32'd70266419);
    Send_IMC_Command(32'd86979380);
    Send_IMC_Command(32'd86912821);
    Send_IMC_Command(32'd87110454);
    Send_IMC_Command(32'd70661431);
    Send_IMC_Command(32'd70529592);
    Send_IMC_Command(32'd70136121);
    Send_IMC_Command(32'd70596922);
    Send_IMC_Command(32'd87372603);
    Send_IMC_Command(32'd70201404);
    Send_IMC_Command(32'd70401085);
    Send_IMC_Command(32'd87175998);
    Send_IMC_Command(32'd86980415);
    Send_IMC_Command(32'd87702336);
    Send_IMC_Command(32'd87111745);
    Send_IMC_Command(32'd87899714);
    Send_IMC_Command(32'd88097347);
    Send_IMC_Command(32'd88031556);
    Send_IMC_Command(32'd88031301);
    Send_IMC_Command(32'd88162886);
    Send_IMC_Command(32'd88359751);
    Send_IMC_Command(32'd71701832);
    Send_IMC_Command(32'd71435849);
    Send_IMC_Command(32'd71373898);
    Send_IMC_Command(32'd71636555);
    Send_IMC_Command(32'd71305292);
    Send_IMC_Command(32'd71241293);
    Send_IMC_Command(32'd71571534);
    Send_IMC_Command(32'd71767887);
    Send_IMC_Command(32'd71502160);
    Send_IMC_Command(32'd71699025);
    Send_IMC_Command(32'd71434322);
    Send_IMC_Command(32'd71370579);
    Send_IMC_Command(32'd71633748);
    Send_IMC_Command(32'd71303509);
    Send_IMC_Command(32'd71241558);
    Send_IMC_Command(32'd71566167);
    Send_IMC_Command(32'd71766104);
    Send_IMC_Command(32'd71500377);
    Send_IMC_Command(32'd89020250);
    Send_IMC_Command(32'd89412955);
    Send_IMC_Command(32'd89151580);
    Send_IMC_Command(32'd88689757);
    Send_IMC_Command(32'd88756830);
    Send_IMC_Command(32'd88624479);
    Send_IMC_Command(32'd88823392);
    Send_IMC_Command(32'd89807713);
    Send_IMC_Command(32'd88887138);
    Send_IMC_Command(32'd89217379);
    Send_IMC_Command(32'd89349732);
    Send_IMC_Command(32'd89808229);
    Send_IMC_Command(32'd88623718);
    Send_IMC_Command(32'd88821095);
    Send_IMC_Command(32'd88823912);
    Send_IMC_Command(32'd89150825);
    Send_IMC_Command(32'd89347946);
    Send_IMC_Command(32'd89414763);
    Send_IMC_Command(32'd89743212);
    Send_IMC_Command(32'd89939309);
    Send_IMC_Command(32'd90071150);
    Send_IMC_Command(32'd89940335);
    Send_IMC_Command(32'd90268272);
    Send_IMC_Command(32'd90136945);
    Send_IMC_Command(32'd90203250);
    Send_IMC_Command(32'd90400115);
    Send_IMC_Command(32'd90467444);
    Send_IMC_Command(32'd90534517);
    Send_IMC_Command(32'd90795638);
    Send_IMC_Command(32'd90664895);
    Send_IMC_Command(32'd91453118);
    Send_IMC_Command(32'd90928573);
    Send_IMC_Command(32'd90599356);
    Send_IMC_Command(32'd91255995);
    Send_IMC_Command(32'd91058618);
    Send_IMC_Command(32'd90730681);
    Send_IMC_Command(32'd90401464);
    Send_IMC_Command(32'd96977920);
    Send_IMC_Command(32'd298238977);
    Send_IMC_Command(32'd298305026);
    Send_IMC_Command(32'd96781059);
    Send_IMC_Command(32'd298041348);
    Send_IMC_Command(32'd96583685);
    Send_IMC_Command(32'd298188806);
    Send_IMC_Command(32'd83952903);
    Send_IMC_Command(32'd297796360);
    Send_IMC_Command(32'd84018185);
    Send_IMC_Command(32'd84018442);
    Send_IMC_Command(32'd84083979);
    Send_IMC_Command(32'd298124044);
    Send_IMC_Command(32'd96911629);
    Send_IMC_Command(32'd298125070);
    Send_IMC_Command(32'd84151567);
    Send_IMC_Command(32'd96667152);
    Send_IMC_Command(32'd298172945);
    Send_IMC_Command(32'd297976082);
    Send_IMC_Command(32'd298173203);
    Send_IMC_Command(32'd96932116);
    Send_IMC_Command(32'd83955989);
    Send_IMC_Command(32'd84742934);
    Send_IMC_Command(32'd84087319);
    Send_IMC_Command(32'd84481816);
    Send_IMC_Command(32'd84480537);
    Send_IMC_Command(32'd84612634);
    Send_IMC_Command(32'd67769627);
    Send_IMC_Command(32'd67110428);
    Send_IMC_Command(32'd85531421);
    Send_IMC_Command(32'd67572766);
    Send_IMC_Command(32'd85859103);
    Send_IMC_Command(32'd67835424);
    Send_IMC_Command(32'd67176481);
    Send_IMC_Command(32'd85598242);
    Send_IMC_Command(32'd68095523);
    Send_IMC_Command(32'd86188068);
    Send_IMC_Command(32'd67311653);
    Send_IMC_Command(32'd68163366);
    Send_IMC_Command(32'd86385959);
    Send_IMC_Command(32'd67242280);
    Send_IMC_Command(32'd86517033);
    Send_IMC_Command(32'd85793834);
    Send_IMC_Command(32'd85918763);
    Send_IMC_Command(32'd86122796);
    Send_IMC_Command(32'd86255917);
    Send_IMC_Command(32'd86648622);
    Send_IMC_Command(32'd86714671);
    Send_IMC_Command(32'd86779696);
    Send_IMC_Command(32'd86838321);
    Send_IMC_Command(32'd87044402);
    Send_IMC_Command(32'd70266419);
    Send_IMC_Command(32'd86979380);
    Send_IMC_Command(32'd86912821);
    Send_IMC_Command(32'd87110454);
    Send_IMC_Command(32'd70661431);
    Send_IMC_Command(32'd70529592);
    Send_IMC_Command(32'd70136121);
    Send_IMC_Command(32'd70596922);
    Send_IMC_Command(32'd87372603);
    Send_IMC_Command(32'd70201404);
    Send_IMC_Command(32'd70401085);
    Send_IMC_Command(32'd87175998);
    Send_IMC_Command(32'd86980415);
    Send_IMC_Command(32'd87702336);
    Send_IMC_Command(32'd87111745);
    Send_IMC_Command(32'd87899714);
    Send_IMC_Command(32'd88097347);
    Send_IMC_Command(32'd88031556);
    Send_IMC_Command(32'd88031301);
    Send_IMC_Command(32'd88162886);
    Send_IMC_Command(32'd88359751);
    Send_IMC_Command(32'd71701832);
    Send_IMC_Command(32'd71435849);
    Send_IMC_Command(32'd71373898);
    Send_IMC_Command(32'd71636555);
    Send_IMC_Command(32'd71305292);
    Send_IMC_Command(32'd71241293);
    Send_IMC_Command(32'd71571534);
    Send_IMC_Command(32'd71767887);
    Send_IMC_Command(32'd71502160);
    Send_IMC_Command(32'd71699025);
    Send_IMC_Command(32'd71434322);
    Send_IMC_Command(32'd71370579);
    Send_IMC_Command(32'd71633748);
    Send_IMC_Command(32'd71303509);
    Send_IMC_Command(32'd71241558);
    Send_IMC_Command(32'd71566167);
    Send_IMC_Command(32'd71766104);
    Send_IMC_Command(32'd71500377);
    Send_IMC_Command(32'd89020250);
    Send_IMC_Command(32'd89412955);
    Send_IMC_Command(32'd89151580);
    Send_IMC_Command(32'd88689757);
    Send_IMC_Command(32'd88756830);
    Send_IMC_Command(32'd88624479);
    Send_IMC_Command(32'd88823392);
    Send_IMC_Command(32'd89807713);
    Send_IMC_Command(32'd88887138);
    Send_IMC_Command(32'd89217379);
    Send_IMC_Command(32'd89349732);
    Send_IMC_Command(32'd89808229);
    Send_IMC_Command(32'd88623718);
    Send_IMC_Command(32'd88821095);
    Send_IMC_Command(32'd88823912);
    Send_IMC_Command(32'd89150825);
    Send_IMC_Command(32'd89347946);
    Send_IMC_Command(32'd89414763);
    Send_IMC_Command(32'd89743212);
    Send_IMC_Command(32'd89939309);
    Send_IMC_Command(32'd90071150);
    Send_IMC_Command(32'd89940335);
    Send_IMC_Command(32'd90268272);
    Send_IMC_Command(32'd90136945);
    Send_IMC_Command(32'd90203250);
    Send_IMC_Command(32'd90400115);
    Send_IMC_Command(32'd90467444);
    Send_IMC_Command(32'd90534517);
    Send_IMC_Command(32'd90795638);
    Send_IMC_Command(32'd90664903);
    Send_IMC_Command(32'd91453126);
    Send_IMC_Command(32'd90928581);
    Send_IMC_Command(32'd90599364);
    Send_IMC_Command(32'd91256003);
    Send_IMC_Command(32'd91058626);
    Send_IMC_Command(32'd90730689);
    Send_IMC_Command(32'd90401472);
    Send_IMC_Command(32'd97504256);
    Send_IMC_Command(32'd298765313);
    Send_IMC_Command(32'd298831362);
    Send_IMC_Command(32'd97307395);
    Send_IMC_Command(32'd298567684);
    Send_IMC_Command(32'd97110021);
    Send_IMC_Command(32'd298713094);
    Send_IMC_Command(32'd83952903);
    Send_IMC_Command(32'd298320648);
    Send_IMC_Command(32'd84018185);
    Send_IMC_Command(32'd84018442);
    Send_IMC_Command(32'd84083979);
    Send_IMC_Command(32'd298648332);
    Send_IMC_Command(32'd97437965);
    Send_IMC_Command(32'd298649358);
    Send_IMC_Command(32'd84151567);
    Send_IMC_Command(32'd97191440);
    Send_IMC_Command(32'd298699281);
    Send_IMC_Command(32'd298502418);
    Send_IMC_Command(32'd298699539);
    Send_IMC_Command(32'd97456404);
    Send_IMC_Command(32'd83955989);
    Send_IMC_Command(32'd84742934);
    Send_IMC_Command(32'd84087319);
    Send_IMC_Command(32'd84481816);
    Send_IMC_Command(32'd84480537);
    Send_IMC_Command(32'd84612634);
    Send_IMC_Command(32'd67769627);
    Send_IMC_Command(32'd67110428);
    Send_IMC_Command(32'd85531421);
    Send_IMC_Command(32'd67572766);
    Send_IMC_Command(32'd85859103);
    Send_IMC_Command(32'd67835424);
    Send_IMC_Command(32'd67176481);
    Send_IMC_Command(32'd85598242);
    Send_IMC_Command(32'd68095523);
    Send_IMC_Command(32'd86188068);
    Send_IMC_Command(32'd67311653);
    Send_IMC_Command(32'd68163366);
    Send_IMC_Command(32'd86385959);
    Send_IMC_Command(32'd67242280);
    Send_IMC_Command(32'd86517033);
    Send_IMC_Command(32'd85793834);
    Send_IMC_Command(32'd85918763);
    Send_IMC_Command(32'd86122796);
    Send_IMC_Command(32'd86255917);
    Send_IMC_Command(32'd86648622);
    Send_IMC_Command(32'd86714671);
    Send_IMC_Command(32'd86779696);
    Send_IMC_Command(32'd86838321);
    Send_IMC_Command(32'd87044402);
    Send_IMC_Command(32'd70266419);
    Send_IMC_Command(32'd86979380);
    Send_IMC_Command(32'd86912821);
    Send_IMC_Command(32'd87110454);
    Send_IMC_Command(32'd70661431);
    Send_IMC_Command(32'd70529592);
    Send_IMC_Command(32'd70136121);
    Send_IMC_Command(32'd70596922);
    Send_IMC_Command(32'd87372603);
    Send_IMC_Command(32'd70201404);
    Send_IMC_Command(32'd70401085);
    Send_IMC_Command(32'd87175998);
    Send_IMC_Command(32'd86980415);
    Send_IMC_Command(32'd87702336);
    Send_IMC_Command(32'd87111745);
    Send_IMC_Command(32'd87899714);
    Send_IMC_Command(32'd88097347);
    Send_IMC_Command(32'd88031556);
    Send_IMC_Command(32'd88031301);
    Send_IMC_Command(32'd88162886);
    Send_IMC_Command(32'd88359751);
    Send_IMC_Command(32'd71701832);
    Send_IMC_Command(32'd71435849);
    Send_IMC_Command(32'd71373898);
    Send_IMC_Command(32'd71636555);
    Send_IMC_Command(32'd71305292);
    Send_IMC_Command(32'd71241293);
    Send_IMC_Command(32'd71571534);
    Send_IMC_Command(32'd71767887);
    Send_IMC_Command(32'd71502160);
    Send_IMC_Command(32'd71699025);
    Send_IMC_Command(32'd71434322);
    Send_IMC_Command(32'd71370579);
    Send_IMC_Command(32'd71633748);
    Send_IMC_Command(32'd71303509);
    Send_IMC_Command(32'd71241558);
    Send_IMC_Command(32'd71566167);
    Send_IMC_Command(32'd71766104);
    Send_IMC_Command(32'd71500377);
    Send_IMC_Command(32'd89020250);
    Send_IMC_Command(32'd89412955);
    Send_IMC_Command(32'd89151580);
    Send_IMC_Command(32'd88689757);
    Send_IMC_Command(32'd88756830);
    Send_IMC_Command(32'd88624479);
    Send_IMC_Command(32'd88823392);
    Send_IMC_Command(32'd89807713);
    Send_IMC_Command(32'd88887138);
    Send_IMC_Command(32'd89217379);
    Send_IMC_Command(32'd89349732);
    Send_IMC_Command(32'd89808229);
    Send_IMC_Command(32'd88623718);
    Send_IMC_Command(32'd88821095);
    Send_IMC_Command(32'd88823912);
    Send_IMC_Command(32'd89150825);
    Send_IMC_Command(32'd89347946);
    Send_IMC_Command(32'd89414763);
    Send_IMC_Command(32'd89743212);
    Send_IMC_Command(32'd89939309);
    Send_IMC_Command(32'd90071150);
    Send_IMC_Command(32'd89940335);
    Send_IMC_Command(32'd90268272);
    Send_IMC_Command(32'd90136945);
    Send_IMC_Command(32'd90203250);
    Send_IMC_Command(32'd90400115);
    Send_IMC_Command(32'd90467444);
    Send_IMC_Command(32'd90534517);
    Send_IMC_Command(32'd90795638);
    Send_IMC_Command(32'd90664911);
    Send_IMC_Command(32'd91453134);
    Send_IMC_Command(32'd90928589);
    Send_IMC_Command(32'd90599372);
    Send_IMC_Command(32'd91256011);
    Send_IMC_Command(32'd91058634);
    Send_IMC_Command(32'd90730697);
    Send_IMC_Command(32'd90401480);
    Send_IMC_Command(32'd98030592);
    Send_IMC_Command(32'd299291649);
    Send_IMC_Command(32'd299357698);
    Send_IMC_Command(32'd97833731);
    Send_IMC_Command(32'd299094020);
    Send_IMC_Command(32'd97636357);
    Send_IMC_Command(32'd299237382);
    Send_IMC_Command(32'd83952903);
    Send_IMC_Command(32'd298844936);
    Send_IMC_Command(32'd84018185);
    Send_IMC_Command(32'd84018442);
    Send_IMC_Command(32'd84083979);
    Send_IMC_Command(32'd299172620);
    Send_IMC_Command(32'd97964301);
    Send_IMC_Command(32'd299173646);
    Send_IMC_Command(32'd84151567);
    Send_IMC_Command(32'd97715728);
    Send_IMC_Command(32'd299225617);
    Send_IMC_Command(32'd299028754);
    Send_IMC_Command(32'd299225875);
    Send_IMC_Command(32'd97980692);
    Send_IMC_Command(32'd83955989);
    Send_IMC_Command(32'd84742934);
    Send_IMC_Command(32'd84087319);
    Send_IMC_Command(32'd84481816);
    Send_IMC_Command(32'd84480537);
    Send_IMC_Command(32'd84612634);
    Send_IMC_Command(32'd67769627);
    Send_IMC_Command(32'd67110428);
    Send_IMC_Command(32'd85531421);
    Send_IMC_Command(32'd67572766);
    Send_IMC_Command(32'd85859103);
    Send_IMC_Command(32'd67835424);
    Send_IMC_Command(32'd67176481);
    Send_IMC_Command(32'd85598242);
    Send_IMC_Command(32'd68095523);
    Send_IMC_Command(32'd86188068);
    Send_IMC_Command(32'd67311653);
    Send_IMC_Command(32'd68163366);
    Send_IMC_Command(32'd86385959);
    Send_IMC_Command(32'd67242280);
    Send_IMC_Command(32'd86517033);
    Send_IMC_Command(32'd85793834);
    Send_IMC_Command(32'd85918763);
    Send_IMC_Command(32'd86122796);
    Send_IMC_Command(32'd86255917);
    Send_IMC_Command(32'd86648622);
    Send_IMC_Command(32'd86714671);
    Send_IMC_Command(32'd86779696);
    Send_IMC_Command(32'd86838321);
    Send_IMC_Command(32'd87044402);
    Send_IMC_Command(32'd70266419);
    Send_IMC_Command(32'd86979380);
    Send_IMC_Command(32'd86912821);
    Send_IMC_Command(32'd87110454);
    Send_IMC_Command(32'd70661431);
    Send_IMC_Command(32'd70529592);
    Send_IMC_Command(32'd70136121);
    Send_IMC_Command(32'd70596922);
    Send_IMC_Command(32'd87372603);
    Send_IMC_Command(32'd70201404);
    Send_IMC_Command(32'd70401085);
    Send_IMC_Command(32'd87175998);
    Send_IMC_Command(32'd86980415);
    Send_IMC_Command(32'd87702336);
    Send_IMC_Command(32'd87111745);
    Send_IMC_Command(32'd87899714);
    Send_IMC_Command(32'd88097347);
    Send_IMC_Command(32'd88031556);
    Send_IMC_Command(32'd88031301);
    Send_IMC_Command(32'd88162886);
    Send_IMC_Command(32'd88359751);
    Send_IMC_Command(32'd71701832);
    Send_IMC_Command(32'd71435849);
    Send_IMC_Command(32'd71373898);
    Send_IMC_Command(32'd71636555);
    Send_IMC_Command(32'd71305292);
    Send_IMC_Command(32'd71241293);
    Send_IMC_Command(32'd71571534);
    Send_IMC_Command(32'd71767887);
    Send_IMC_Command(32'd71502160);
    Send_IMC_Command(32'd71699025);
    Send_IMC_Command(32'd71434322);
    Send_IMC_Command(32'd71370579);
    Send_IMC_Command(32'd71633748);
    Send_IMC_Command(32'd71303509);
    Send_IMC_Command(32'd71241558);
    Send_IMC_Command(32'd71566167);
    Send_IMC_Command(32'd71766104);
    Send_IMC_Command(32'd71500377);
    Send_IMC_Command(32'd89020250);
    Send_IMC_Command(32'd89412955);
    Send_IMC_Command(32'd89151580);
    Send_IMC_Command(32'd88689757);
    Send_IMC_Command(32'd88756830);
    Send_IMC_Command(32'd88624479);
    Send_IMC_Command(32'd88823392);
    Send_IMC_Command(32'd89807713);
    Send_IMC_Command(32'd88887138);
    Send_IMC_Command(32'd89217379);
    Send_IMC_Command(32'd89349732);
    Send_IMC_Command(32'd89808229);
    Send_IMC_Command(32'd88623718);
    Send_IMC_Command(32'd88821095);
    Send_IMC_Command(32'd88823912);
    Send_IMC_Command(32'd89150825);
    Send_IMC_Command(32'd89347946);
    Send_IMC_Command(32'd89414763);
    Send_IMC_Command(32'd89743212);
    Send_IMC_Command(32'd89939309);
    Send_IMC_Command(32'd90071150);
    Send_IMC_Command(32'd89940335);
    Send_IMC_Command(32'd90268272);
    Send_IMC_Command(32'd90136945);
    Send_IMC_Command(32'd90203250);
    Send_IMC_Command(32'd90400115);
    Send_IMC_Command(32'd90467444);
    Send_IMC_Command(32'd90534517);
    Send_IMC_Command(32'd90795638);
    Send_IMC_Command(32'd90664919);
    Send_IMC_Command(32'd91453142);
    Send_IMC_Command(32'd90928597);
    Send_IMC_Command(32'd90599380);
    Send_IMC_Command(32'd91256019);
    Send_IMC_Command(32'd91058642);
    Send_IMC_Command(32'd90730705);
    Send_IMC_Command(32'd90401488);
    Send_IMC_Command(32'd98556928);
    Send_IMC_Command(32'd299817985);
    Send_IMC_Command(32'd299884034);
    Send_IMC_Command(32'd98360067);
    Send_IMC_Command(32'd299620356);
    Send_IMC_Command(32'd98162693);
    Send_IMC_Command(32'd299761670);
    Send_IMC_Command(32'd83952903);
    Send_IMC_Command(32'd299369224);
    Send_IMC_Command(32'd84018185);
    Send_IMC_Command(32'd84018442);
    Send_IMC_Command(32'd84083979);
    Send_IMC_Command(32'd299696908);
    Send_IMC_Command(32'd98490637);
    Send_IMC_Command(32'd299697934);
    Send_IMC_Command(32'd84151567);
    Send_IMC_Command(32'd98240016);
    Send_IMC_Command(32'd299751953);
    Send_IMC_Command(32'd299555090);
    Send_IMC_Command(32'd299752211);
    Send_IMC_Command(32'd98504980);
    Send_IMC_Command(32'd83955989);
    Send_IMC_Command(32'd84742934);
    Send_IMC_Command(32'd84087319);
    Send_IMC_Command(32'd84481816);
    Send_IMC_Command(32'd84480537);
    Send_IMC_Command(32'd84612634);
    Send_IMC_Command(32'd67769627);
    Send_IMC_Command(32'd67110428);
    Send_IMC_Command(32'd85531421);
    Send_IMC_Command(32'd67572766);
    Send_IMC_Command(32'd85859103);
    Send_IMC_Command(32'd67835424);
    Send_IMC_Command(32'd67176481);
    Send_IMC_Command(32'd85598242);
    Send_IMC_Command(32'd68095523);
    Send_IMC_Command(32'd86188068);
    Send_IMC_Command(32'd67311653);
    Send_IMC_Command(32'd68163366);
    Send_IMC_Command(32'd86385959);
    Send_IMC_Command(32'd67242280);
    Send_IMC_Command(32'd86517033);
    Send_IMC_Command(32'd85793834);
    Send_IMC_Command(32'd85918763);
    Send_IMC_Command(32'd86122796);
    Send_IMC_Command(32'd86255917);
    Send_IMC_Command(32'd86648622);
    Send_IMC_Command(32'd86714671);
    Send_IMC_Command(32'd86779696);
    Send_IMC_Command(32'd86838321);
    Send_IMC_Command(32'd87044402);
    Send_IMC_Command(32'd70266419);
    Send_IMC_Command(32'd86979380);
    Send_IMC_Command(32'd86912821);
    Send_IMC_Command(32'd87110454);
    Send_IMC_Command(32'd70661431);
    Send_IMC_Command(32'd70529592);
    Send_IMC_Command(32'd70136121);
    Send_IMC_Command(32'd70596922);
    Send_IMC_Command(32'd87372603);
    Send_IMC_Command(32'd70201404);
    Send_IMC_Command(32'd70401085);
    Send_IMC_Command(32'd87175998);
    Send_IMC_Command(32'd86980415);
    Send_IMC_Command(32'd87702336);
    Send_IMC_Command(32'd87111745);
    Send_IMC_Command(32'd87899714);
    Send_IMC_Command(32'd88097347);
    Send_IMC_Command(32'd88031556);
    Send_IMC_Command(32'd88031301);
    Send_IMC_Command(32'd88162886);
    Send_IMC_Command(32'd88359751);
    Send_IMC_Command(32'd71701832);
    Send_IMC_Command(32'd71435849);
    Send_IMC_Command(32'd71373898);
    Send_IMC_Command(32'd71636555);
    Send_IMC_Command(32'd71305292);
    Send_IMC_Command(32'd71241293);
    Send_IMC_Command(32'd71571534);
    Send_IMC_Command(32'd71767887);
    Send_IMC_Command(32'd71502160);
    Send_IMC_Command(32'd71699025);
    Send_IMC_Command(32'd71434322);
    Send_IMC_Command(32'd71370579);
    Send_IMC_Command(32'd71633748);
    Send_IMC_Command(32'd71303509);
    Send_IMC_Command(32'd71241558);
    Send_IMC_Command(32'd71566167);
    Send_IMC_Command(32'd71766104);
    Send_IMC_Command(32'd71500377);
    Send_IMC_Command(32'd89020250);
    Send_IMC_Command(32'd89412955);
    Send_IMC_Command(32'd89151580);
    Send_IMC_Command(32'd88689757);
    Send_IMC_Command(32'd88756830);
    Send_IMC_Command(32'd88624479);
    Send_IMC_Command(32'd88823392);
    Send_IMC_Command(32'd89807713);
    Send_IMC_Command(32'd88887138);
    Send_IMC_Command(32'd89217379);
    Send_IMC_Command(32'd89349732);
    Send_IMC_Command(32'd89808229);
    Send_IMC_Command(32'd88623718);
    Send_IMC_Command(32'd88821095);
    Send_IMC_Command(32'd88823912);
    Send_IMC_Command(32'd89150825);
    Send_IMC_Command(32'd89347946);
    Send_IMC_Command(32'd89414763);
    Send_IMC_Command(32'd89743212);
    Send_IMC_Command(32'd89939309);
    Send_IMC_Command(32'd90071150);
    Send_IMC_Command(32'd89940335);
    Send_IMC_Command(32'd90268272);
    Send_IMC_Command(32'd90136945);
    Send_IMC_Command(32'd90203250);
    Send_IMC_Command(32'd90400115);
    Send_IMC_Command(32'd90467444);
    Send_IMC_Command(32'd90534517);
    Send_IMC_Command(32'd90795638);
    Send_IMC_Command(32'd90664927);
    Send_IMC_Command(32'd91453150);
    Send_IMC_Command(32'd90928605);
    Send_IMC_Command(32'd90599388);
    Send_IMC_Command(32'd91256027);
    Send_IMC_Command(32'd91058650);
    Send_IMC_Command(32'd90730713);
    Send_IMC_Command(32'd90401496);
    Send_IMC_Command(32'd99083264);
    Send_IMC_Command(32'd300344321);
    Send_IMC_Command(32'd300410370);
    Send_IMC_Command(32'd98886403);
    Send_IMC_Command(32'd300146692);
    Send_IMC_Command(32'd98689029);
    Send_IMC_Command(32'd300285958);
    Send_IMC_Command(32'd83952903);
    Send_IMC_Command(32'd299893512);
    Send_IMC_Command(32'd84018185);
    Send_IMC_Command(32'd84018442);
    Send_IMC_Command(32'd84083979);
    Send_IMC_Command(32'd300221196);
    Send_IMC_Command(32'd99016973);
    Send_IMC_Command(32'd300222222);
    Send_IMC_Command(32'd84151567);
    Send_IMC_Command(32'd98764304);
    Send_IMC_Command(32'd300278289);
    Send_IMC_Command(32'd300081426);
    Send_IMC_Command(32'd300278547);
    Send_IMC_Command(32'd99029268);
    Send_IMC_Command(32'd83955989);
    Send_IMC_Command(32'd84742934);
    Send_IMC_Command(32'd84087319);
    Send_IMC_Command(32'd84481816);
    Send_IMC_Command(32'd84480537);
    Send_IMC_Command(32'd84612634);
    Send_IMC_Command(32'd67769627);
    Send_IMC_Command(32'd67110428);
    Send_IMC_Command(32'd85531421);
    Send_IMC_Command(32'd67572766);
    Send_IMC_Command(32'd85859103);
    Send_IMC_Command(32'd67835424);
    Send_IMC_Command(32'd67176481);
    Send_IMC_Command(32'd85598242);
    Send_IMC_Command(32'd68095523);
    Send_IMC_Command(32'd86188068);
    Send_IMC_Command(32'd67311653);
    Send_IMC_Command(32'd68163366);
    Send_IMC_Command(32'd86385959);
    Send_IMC_Command(32'd67242280);
    Send_IMC_Command(32'd86517033);
    Send_IMC_Command(32'd85793834);
    Send_IMC_Command(32'd85918763);
    Send_IMC_Command(32'd86122796);
    Send_IMC_Command(32'd86255917);
    Send_IMC_Command(32'd86648622);
    Send_IMC_Command(32'd86714671);
    Send_IMC_Command(32'd86779696);
    Send_IMC_Command(32'd86838321);
    Send_IMC_Command(32'd87044402);
    Send_IMC_Command(32'd70266419);
    Send_IMC_Command(32'd86979380);
    Send_IMC_Command(32'd86912821);
    Send_IMC_Command(32'd87110454);
    Send_IMC_Command(32'd70661431);
    Send_IMC_Command(32'd70529592);
    Send_IMC_Command(32'd70136121);
    Send_IMC_Command(32'd70596922);
    Send_IMC_Command(32'd87372603);
    Send_IMC_Command(32'd70201404);
    Send_IMC_Command(32'd70401085);
    Send_IMC_Command(32'd87175998);
    Send_IMC_Command(32'd86980415);
    Send_IMC_Command(32'd87702336);
    Send_IMC_Command(32'd87111745);
    Send_IMC_Command(32'd87899714);
    Send_IMC_Command(32'd88097347);
    Send_IMC_Command(32'd88031556);
    Send_IMC_Command(32'd88031301);
    Send_IMC_Command(32'd88162886);
    Send_IMC_Command(32'd88359751);
    Send_IMC_Command(32'd71701832);
    Send_IMC_Command(32'd71435849);
    Send_IMC_Command(32'd71373898);
    Send_IMC_Command(32'd71636555);
    Send_IMC_Command(32'd71305292);
    Send_IMC_Command(32'd71241293);
    Send_IMC_Command(32'd71571534);
    Send_IMC_Command(32'd71767887);
    Send_IMC_Command(32'd71502160);
    Send_IMC_Command(32'd71699025);
    Send_IMC_Command(32'd71434322);
    Send_IMC_Command(32'd71370579);
    Send_IMC_Command(32'd71633748);
    Send_IMC_Command(32'd71303509);
    Send_IMC_Command(32'd71241558);
    Send_IMC_Command(32'd71566167);
    Send_IMC_Command(32'd71766104);
    Send_IMC_Command(32'd71500377);
    Send_IMC_Command(32'd89020250);
    Send_IMC_Command(32'd89412955);
    Send_IMC_Command(32'd89151580);
    Send_IMC_Command(32'd88689757);
    Send_IMC_Command(32'd88756830);
    Send_IMC_Command(32'd88624479);
    Send_IMC_Command(32'd88823392);
    Send_IMC_Command(32'd89807713);
    Send_IMC_Command(32'd88887138);
    Send_IMC_Command(32'd89217379);
    Send_IMC_Command(32'd89349732);
    Send_IMC_Command(32'd89808229);
    Send_IMC_Command(32'd88623718);
    Send_IMC_Command(32'd88821095);
    Send_IMC_Command(32'd88823912);
    Send_IMC_Command(32'd89150825);
    Send_IMC_Command(32'd89347946);
    Send_IMC_Command(32'd89414763);
    Send_IMC_Command(32'd89743212);
    Send_IMC_Command(32'd89939309);
    Send_IMC_Command(32'd90071150);
    Send_IMC_Command(32'd89940335);
    Send_IMC_Command(32'd90268272);
    Send_IMC_Command(32'd90136945);
    Send_IMC_Command(32'd90203250);
    Send_IMC_Command(32'd90400115);
    Send_IMC_Command(32'd90467444);
    Send_IMC_Command(32'd90534517);
    Send_IMC_Command(32'd90795638);
    Send_IMC_Command(32'd90664935);
    Send_IMC_Command(32'd91453158);
    Send_IMC_Command(32'd90928613);
    Send_IMC_Command(32'd90599396);
    Send_IMC_Command(32'd91256035);
    Send_IMC_Command(32'd91058658);
    Send_IMC_Command(32'd90730721);
    Send_IMC_Command(32'd90401504);
    Send_IMC_Command(32'd99609600);
    Send_IMC_Command(32'd300870657);
    Send_IMC_Command(32'd300936706);
    Send_IMC_Command(32'd99412739);
    Send_IMC_Command(32'd300673028);
    Send_IMC_Command(32'd99215365);
    Send_IMC_Command(32'd300810246);
    Send_IMC_Command(32'd83952903);
    Send_IMC_Command(32'd300417800);
    Send_IMC_Command(32'd84018185);
    Send_IMC_Command(32'd84018442);
    Send_IMC_Command(32'd84083979);
    Send_IMC_Command(32'd300745484);
    Send_IMC_Command(32'd99543309);
    Send_IMC_Command(32'd300746510);
    Send_IMC_Command(32'd84151567);
    Send_IMC_Command(32'd99288592);
    Send_IMC_Command(32'd300804625);
    Send_IMC_Command(32'd300607762);
    Send_IMC_Command(32'd300804883);
    Send_IMC_Command(32'd99553556);
    Send_IMC_Command(32'd83955989);
    Send_IMC_Command(32'd84742934);
    Send_IMC_Command(32'd84087319);
    Send_IMC_Command(32'd84481816);
    Send_IMC_Command(32'd84480537);
    Send_IMC_Command(32'd84612634);
    Send_IMC_Command(32'd67769627);
    Send_IMC_Command(32'd67110428);
    Send_IMC_Command(32'd85531421);
    Send_IMC_Command(32'd67572766);
    Send_IMC_Command(32'd85859103);
    Send_IMC_Command(32'd67835424);
    Send_IMC_Command(32'd67176481);
    Send_IMC_Command(32'd85598242);
    Send_IMC_Command(32'd68095523);
    Send_IMC_Command(32'd86188068);
    Send_IMC_Command(32'd67311653);
    Send_IMC_Command(32'd68163366);
    Send_IMC_Command(32'd86385959);
    Send_IMC_Command(32'd67242280);
    Send_IMC_Command(32'd86517033);
    Send_IMC_Command(32'd85793834);
    Send_IMC_Command(32'd85918763);
    Send_IMC_Command(32'd86122796);
    Send_IMC_Command(32'd86255917);
    Send_IMC_Command(32'd86648622);
    Send_IMC_Command(32'd86714671);
    Send_IMC_Command(32'd86779696);
    Send_IMC_Command(32'd86838321);
    Send_IMC_Command(32'd87044402);
    Send_IMC_Command(32'd70266419);
    Send_IMC_Command(32'd86979380);
    Send_IMC_Command(32'd86912821);
    Send_IMC_Command(32'd87110454);
    Send_IMC_Command(32'd70661431);
    Send_IMC_Command(32'd70529592);
    Send_IMC_Command(32'd70136121);
    Send_IMC_Command(32'd70596922);
    Send_IMC_Command(32'd87372603);
    Send_IMC_Command(32'd70201404);
    Send_IMC_Command(32'd70401085);
    Send_IMC_Command(32'd87175998);
    Send_IMC_Command(32'd86980415);
    Send_IMC_Command(32'd87702336);
    Send_IMC_Command(32'd87111745);
    Send_IMC_Command(32'd87899714);
    Send_IMC_Command(32'd88097347);
    Send_IMC_Command(32'd88031556);
    Send_IMC_Command(32'd88031301);
    Send_IMC_Command(32'd88162886);
    Send_IMC_Command(32'd88359751);
    Send_IMC_Command(32'd71701832);
    Send_IMC_Command(32'd71435849);
    Send_IMC_Command(32'd71373898);
    Send_IMC_Command(32'd71636555);
    Send_IMC_Command(32'd71305292);
    Send_IMC_Command(32'd71241293);
    Send_IMC_Command(32'd71571534);
    Send_IMC_Command(32'd71767887);
    Send_IMC_Command(32'd71502160);
    Send_IMC_Command(32'd71699025);
    Send_IMC_Command(32'd71434322);
    Send_IMC_Command(32'd71370579);
    Send_IMC_Command(32'd71633748);
    Send_IMC_Command(32'd71303509);
    Send_IMC_Command(32'd71241558);
    Send_IMC_Command(32'd71566167);
    Send_IMC_Command(32'd71766104);
    Send_IMC_Command(32'd71500377);
    Send_IMC_Command(32'd89020250);
    Send_IMC_Command(32'd89412955);
    Send_IMC_Command(32'd89151580);
    Send_IMC_Command(32'd88689757);
    Send_IMC_Command(32'd88756830);
    Send_IMC_Command(32'd88624479);
    Send_IMC_Command(32'd88823392);
    Send_IMC_Command(32'd89807713);
    Send_IMC_Command(32'd88887138);
    Send_IMC_Command(32'd89217379);
    Send_IMC_Command(32'd89349732);
    Send_IMC_Command(32'd89808229);
    Send_IMC_Command(32'd88623718);
    Send_IMC_Command(32'd88821095);
    Send_IMC_Command(32'd88823912);
    Send_IMC_Command(32'd89150825);
    Send_IMC_Command(32'd89347946);
    Send_IMC_Command(32'd89414763);
    Send_IMC_Command(32'd89743212);
    Send_IMC_Command(32'd89939309);
    Send_IMC_Command(32'd90071150);
    Send_IMC_Command(32'd89940335);
    Send_IMC_Command(32'd90268272);
    Send_IMC_Command(32'd90136945);
    Send_IMC_Command(32'd90203250);
    Send_IMC_Command(32'd90400115);
    Send_IMC_Command(32'd90467444);
    Send_IMC_Command(32'd90534517);
    Send_IMC_Command(32'd90795638);
    Send_IMC_Command(32'd90664943);
    Send_IMC_Command(32'd91453166);
    Send_IMC_Command(32'd90928621);
    Send_IMC_Command(32'd90599404);
    Send_IMC_Command(32'd91256043);
    Send_IMC_Command(32'd91058666);
    Send_IMC_Command(32'd90730729);
    Send_IMC_Command(32'd90401512);
    Send_IMC_Command(32'd100135936);
    Send_IMC_Command(32'd301396993);
    Send_IMC_Command(32'd301463042);
    Send_IMC_Command(32'd99939075);
    Send_IMC_Command(32'd301199364);
    Send_IMC_Command(32'd99741701);
    Send_IMC_Command(32'd301334534);
    Send_IMC_Command(32'd83952903);
    Send_IMC_Command(32'd300942088);
    Send_IMC_Command(32'd84018185);
    Send_IMC_Command(32'd84018442);
    Send_IMC_Command(32'd84083979);
    Send_IMC_Command(32'd301269772);
    Send_IMC_Command(32'd100069645);
    Send_IMC_Command(32'd301270798);
    Send_IMC_Command(32'd84151567);
    Send_IMC_Command(32'd99812880);
    Send_IMC_Command(32'd301330961);
    Send_IMC_Command(32'd301134098);
    Send_IMC_Command(32'd301331219);
    Send_IMC_Command(32'd100077844);
    Send_IMC_Command(32'd83955989);
    Send_IMC_Command(32'd84742934);
    Send_IMC_Command(32'd84087319);
    Send_IMC_Command(32'd84481816);
    Send_IMC_Command(32'd84480537);
    Send_IMC_Command(32'd84612634);
    Send_IMC_Command(32'd67769627);
    Send_IMC_Command(32'd67110428);
    Send_IMC_Command(32'd85531421);
    Send_IMC_Command(32'd67572766);
    Send_IMC_Command(32'd85859103);
    Send_IMC_Command(32'd67835424);
    Send_IMC_Command(32'd67176481);
    Send_IMC_Command(32'd85598242);
    Send_IMC_Command(32'd68095523);
    Send_IMC_Command(32'd86188068);
    Send_IMC_Command(32'd67311653);
    Send_IMC_Command(32'd68163366);
    Send_IMC_Command(32'd86385959);
    Send_IMC_Command(32'd67242280);
    Send_IMC_Command(32'd86517033);
    Send_IMC_Command(32'd85793834);
    Send_IMC_Command(32'd85918763);
    Send_IMC_Command(32'd86122796);
    Send_IMC_Command(32'd86255917);
    Send_IMC_Command(32'd86648622);
    Send_IMC_Command(32'd86714671);
    Send_IMC_Command(32'd86779696);
    Send_IMC_Command(32'd86838321);
    Send_IMC_Command(32'd87044402);
    Send_IMC_Command(32'd70266419);
    Send_IMC_Command(32'd86979380);
    Send_IMC_Command(32'd86912821);
    Send_IMC_Command(32'd87110454);
    Send_IMC_Command(32'd70661431);
    Send_IMC_Command(32'd70529592);
    Send_IMC_Command(32'd70136121);
    Send_IMC_Command(32'd70596922);
    Send_IMC_Command(32'd87372603);
    Send_IMC_Command(32'd70201404);
    Send_IMC_Command(32'd70401085);
    Send_IMC_Command(32'd87175998);
    Send_IMC_Command(32'd86980415);
    Send_IMC_Command(32'd87702336);
    Send_IMC_Command(32'd87111745);
    Send_IMC_Command(32'd87899714);
    Send_IMC_Command(32'd88097347);
    Send_IMC_Command(32'd88031556);
    Send_IMC_Command(32'd88031301);
    Send_IMC_Command(32'd88162886);
    Send_IMC_Command(32'd88359751);
    Send_IMC_Command(32'd71701832);
    Send_IMC_Command(32'd71435849);
    Send_IMC_Command(32'd71373898);
    Send_IMC_Command(32'd71636555);
    Send_IMC_Command(32'd71305292);
    Send_IMC_Command(32'd71241293);
    Send_IMC_Command(32'd71571534);
    Send_IMC_Command(32'd71767887);
    Send_IMC_Command(32'd71502160);
    Send_IMC_Command(32'd71699025);
    Send_IMC_Command(32'd71434322);
    Send_IMC_Command(32'd71370579);
    Send_IMC_Command(32'd71633748);
    Send_IMC_Command(32'd71303509);
    Send_IMC_Command(32'd71241558);
    Send_IMC_Command(32'd71566167);
    Send_IMC_Command(32'd71766104);
    Send_IMC_Command(32'd71500377);
    Send_IMC_Command(32'd89020250);
    Send_IMC_Command(32'd89412955);
    Send_IMC_Command(32'd89151580);
    Send_IMC_Command(32'd88689757);
    Send_IMC_Command(32'd88756830);
    Send_IMC_Command(32'd88624479);
    Send_IMC_Command(32'd88823392);
    Send_IMC_Command(32'd89807713);
    Send_IMC_Command(32'd88887138);
    Send_IMC_Command(32'd89217379);
    Send_IMC_Command(32'd89349732);
    Send_IMC_Command(32'd89808229);
    Send_IMC_Command(32'd88623718);
    Send_IMC_Command(32'd88821095);
    Send_IMC_Command(32'd88823912);
    Send_IMC_Command(32'd89150825);
    Send_IMC_Command(32'd89347946);
    Send_IMC_Command(32'd89414763);
    Send_IMC_Command(32'd89743212);
    Send_IMC_Command(32'd89939309);
    Send_IMC_Command(32'd90071150);
    Send_IMC_Command(32'd89940335);
    Send_IMC_Command(32'd90268272);
    Send_IMC_Command(32'd90136945);
    Send_IMC_Command(32'd90203250);
    Send_IMC_Command(32'd90400115);
    Send_IMC_Command(32'd90467444);
    Send_IMC_Command(32'd90534517);
    Send_IMC_Command(32'd90795638);
    Send_IMC_Command(32'd90664951);
    Send_IMC_Command(32'd91453174);
    Send_IMC_Command(32'd90928629);
    Send_IMC_Command(32'd90599412);
    Send_IMC_Command(32'd91256051);
    Send_IMC_Command(32'd91058674);
    Send_IMC_Command(32'd90730737);
    Send_IMC_Command(32'd90401520);
    Send_IMC_Command(32'd100662272);
    Send_IMC_Command(32'd301923329);
    Send_IMC_Command(32'd301989378);
    Send_IMC_Command(32'd100465411);
    Send_IMC_Command(32'd301725700);
    Send_IMC_Command(32'd100268037);
    Send_IMC_Command(32'd301858822);
    Send_IMC_Command(32'd83952903);
    Send_IMC_Command(32'd301466376);
    Send_IMC_Command(32'd84018185);
    Send_IMC_Command(32'd84018442);
    Send_IMC_Command(32'd84083979);
    Send_IMC_Command(32'd301794060);
    Send_IMC_Command(32'd100595981);
    Send_IMC_Command(32'd301795086);
    Send_IMC_Command(32'd84151567);
    Send_IMC_Command(32'd100337168);
    Send_IMC_Command(32'd301857297);
    Send_IMC_Command(32'd301660434);
    Send_IMC_Command(32'd301857555);
    Send_IMC_Command(32'd100602132);
    Send_IMC_Command(32'd83955989);
    Send_IMC_Command(32'd84742934);
    Send_IMC_Command(32'd84087319);
    Send_IMC_Command(32'd84481816);
    Send_IMC_Command(32'd84480537);
    Send_IMC_Command(32'd84612634);
    Send_IMC_Command(32'd67769627);
    Send_IMC_Command(32'd67110428);
    Send_IMC_Command(32'd85531421);
    Send_IMC_Command(32'd67572766);
    Send_IMC_Command(32'd85859103);
    Send_IMC_Command(32'd67835424);
    Send_IMC_Command(32'd67176481);
    Send_IMC_Command(32'd85598242);
    Send_IMC_Command(32'd68095523);
    Send_IMC_Command(32'd86188068);
    Send_IMC_Command(32'd67311653);
    Send_IMC_Command(32'd68163366);
    Send_IMC_Command(32'd86385959);
    Send_IMC_Command(32'd67242280);
    Send_IMC_Command(32'd86517033);
    Send_IMC_Command(32'd85793834);
    Send_IMC_Command(32'd85918763);
    Send_IMC_Command(32'd86122796);
    Send_IMC_Command(32'd86255917);
    Send_IMC_Command(32'd86648622);
    Send_IMC_Command(32'd86714671);
    Send_IMC_Command(32'd86779696);
    Send_IMC_Command(32'd86838321);
    Send_IMC_Command(32'd87044402);
    Send_IMC_Command(32'd70266419);
    Send_IMC_Command(32'd86979380);
    Send_IMC_Command(32'd86912821);
    Send_IMC_Command(32'd87110454);
    Send_IMC_Command(32'd70661431);
    Send_IMC_Command(32'd70529592);
    Send_IMC_Command(32'd70136121);
    Send_IMC_Command(32'd70596922);
    Send_IMC_Command(32'd87372603);
    Send_IMC_Command(32'd70201404);
    Send_IMC_Command(32'd70401085);
    Send_IMC_Command(32'd87175998);
    Send_IMC_Command(32'd86980415);
    Send_IMC_Command(32'd87702336);
    Send_IMC_Command(32'd87111745);
    Send_IMC_Command(32'd87899714);
    Send_IMC_Command(32'd88097347);
    Send_IMC_Command(32'd88031556);
    Send_IMC_Command(32'd88031301);
    Send_IMC_Command(32'd88162886);
    Send_IMC_Command(32'd88359751);
    Send_IMC_Command(32'd71701832);
    Send_IMC_Command(32'd71435849);
    Send_IMC_Command(32'd71373898);
    Send_IMC_Command(32'd71636555);
    Send_IMC_Command(32'd71305292);
    Send_IMC_Command(32'd71241293);
    Send_IMC_Command(32'd71571534);
    Send_IMC_Command(32'd71767887);
    Send_IMC_Command(32'd71502160);
    Send_IMC_Command(32'd71699025);
    Send_IMC_Command(32'd71434322);
    Send_IMC_Command(32'd71370579);
    Send_IMC_Command(32'd71633748);
    Send_IMC_Command(32'd71303509);
    Send_IMC_Command(32'd71241558);
    Send_IMC_Command(32'd71566167);
    Send_IMC_Command(32'd71766104);
    Send_IMC_Command(32'd71500377);
    Send_IMC_Command(32'd89020250);
    Send_IMC_Command(32'd89412955);
    Send_IMC_Command(32'd89151580);
    Send_IMC_Command(32'd88689757);
    Send_IMC_Command(32'd88756830);
    Send_IMC_Command(32'd88624479);
    Send_IMC_Command(32'd88823392);
    Send_IMC_Command(32'd89807713);
    Send_IMC_Command(32'd88887138);
    Send_IMC_Command(32'd89217379);
    Send_IMC_Command(32'd89349732);
    Send_IMC_Command(32'd89808229);
    Send_IMC_Command(32'd88623718);
    Send_IMC_Command(32'd88821095);
    Send_IMC_Command(32'd88823912);
    Send_IMC_Command(32'd89150825);
    Send_IMC_Command(32'd89347946);
    Send_IMC_Command(32'd89414763);
    Send_IMC_Command(32'd89743212);
    Send_IMC_Command(32'd89939309);
    Send_IMC_Command(32'd90071150);
    Send_IMC_Command(32'd89940335);
    Send_IMC_Command(32'd90268272);
    Send_IMC_Command(32'd90136945);
    Send_IMC_Command(32'd90203250);
    Send_IMC_Command(32'd90400115);
    Send_IMC_Command(32'd90467444);
    Send_IMC_Command(32'd90534517);
    Send_IMC_Command(32'd90795638);
    Send_IMC_Command(32'd90664959);
    Send_IMC_Command(32'd91453182);
    Send_IMC_Command(32'd90928637);
    Send_IMC_Command(32'd90599420);
    Send_IMC_Command(32'd91256059);
    Send_IMC_Command(32'd91058682);
    Send_IMC_Command(32'd90730745);
    Send_IMC_Command(32'd90401528);

endtask


task AES_Inv_MC();

    Send_IMC_Command(32'd83888264);
    Send_IMC_Command(32'd84940937);
    Send_IMC_Command(32'd83954058);
    Send_IMC_Command(32'd85006731);
    Send_IMC_Command(32'd84019852);
    Send_IMC_Command(32'd85072525);
    Send_IMC_Command(32'd84085646);
    Send_IMC_Command(32'd85138319);
    Send_IMC_Command(32'd84151440);
    Send_IMC_Command(32'd85204113);
    Send_IMC_Command(32'd84217234);
    Send_IMC_Command(32'd85269907);
    Send_IMC_Command(32'd84283028);
    Send_IMC_Command(32'd85335701);
    Send_IMC_Command(32'd85401494);
    Send_IMC_Command(32'd84348823);
    Send_IMC_Command(32'd84445592);
    Send_IMC_Command(32'd93821056);
    Send_IMC_Command(32'd84350873);
    Send_IMC_Command(32'd85493914);
    Send_IMC_Command(32'd93756112);
    Send_IMC_Command(32'd92917915);
    Send_IMC_Command(32'd93953016);
    Send_IMC_Command(32'd85694108);
    Send_IMC_Command(32'd92831901);
    Send_IMC_Command(32'd93953448);
    Send_IMC_Command(32'd93166750);
    Send_IMC_Command(32'd93232851);
    Send_IMC_Command(32'd84645791);
    Send_IMC_Command(32'd93298592);
    Send_IMC_Command(32'd93102211);
    Send_IMC_Command(32'd84021921);
    Send_IMC_Command(32'd93954466);
    Send_IMC_Command(32'd93429667);
    Send_IMC_Command(32'd93363364);
    Send_IMC_Command(32'd84576933);
    Send_IMC_Command(32'd93169026);
    Send_IMC_Command(32'd85625766);
    Send_IMC_Command(32'd93103826);
    Send_IMC_Command(32'd84482471);
    Send_IMC_Command(32'd94480304);
    Send_IMC_Command(32'd94810282);
    Send_IMC_Command(32'd94744826);
    Send_IMC_Command(32'd83991217);
    Send_IMC_Command(32'd85889970);
    Send_IMC_Command(32'd93631190);
    Send_IMC_Command(32'd84841907);
    Send_IMC_Command(32'd93500294);
    Send_IMC_Command(32'd84219316);
    Send_IMC_Command(32'd85891509);
    Send_IMC_Command(32'd85039286);
    Send_IMC_Command(32'd84775095);
    Send_IMC_Command(32'd93566853);
    Send_IMC_Command(32'd84718776);
    Send_IMC_Command(32'd85823929);
    Send_IMC_Command(32'd93501909);
    Send_IMC_Command(32'd85768378);
    Send_IMC_Command(32'd96058029);
    Send_IMC_Command(32'd95927037);
    Send_IMC_Command(32'd84907195);
    Send_IMC_Command(32'd93764487);
    Send_IMC_Command(32'd84850108);
    Send_IMC_Command(32'd96189695);
    Send_IMC_Command(32'd85956029);
    Send_IMC_Command(32'd96255407);
    Send_IMC_Command(32'd93830615);
    Send_IMC_Command(32'd93631678);
    Send_IMC_Command(32'd92716718);
    Send_IMC_Command(32'd94876095);
    Send_IMC_Command(32'd94093265);
    Send_IMC_Command(32'd93225920);
    Send_IMC_Command(32'd94552235);
    Send_IMC_Command(32'd92976833);
    Send_IMC_Command(32'd100188665);
    Send_IMC_Command(32'd93311938);
    Send_IMC_Command(32'd94552827);
    Send_IMC_Command(32'd85376707);
    Send_IMC_Command(32'd93570046);
    Send_IMC_Command(32'd85173444);
    Send_IMC_Command(32'd85771476);
    Send_IMC_Command(32'd84124613);
    Send_IMC_Command(32'd84723076);
    Send_IMC_Command(32'd93041094);
    Send_IMC_Command(32'd94946985);
    Send_IMC_Command(32'd94218183);
    Send_IMC_Command(32'd95864705);
    Send_IMC_Command(32'd84187592);
    Send_IMC_Command(32'd85182665);
    Send_IMC_Command(32'd94620076);
    Send_IMC_Command(32'd84124874);
    Send_IMC_Command(32'd93965003);
    Send_IMC_Command(32'd85249020);
    Send_IMC_Command(32'd92317832);
    Send_IMC_Command(32'd97581193);
    Send_IMC_Command(32'd92383626);
    Send_IMC_Command(32'd97646987);
    Send_IMC_Command(32'd92449420);
    Send_IMC_Command(32'd97712781);
    Send_IMC_Command(32'd92515214);
    Send_IMC_Command(32'd97778575);
    Send_IMC_Command(32'd92581008);
    Send_IMC_Command(32'd97844369);
    Send_IMC_Command(32'd92646802);
    Send_IMC_Command(32'd97910163);
    Send_IMC_Command(32'd92712596);
    Send_IMC_Command(32'd97975957);
    Send_IMC_Command(32'd98041750);
    Send_IMC_Command(32'd92778391);
    Send_IMC_Command(32'd94931352);
    Send_IMC_Command(32'd93820928);
    Send_IMC_Command(32'd92788633);
    Send_IMC_Command(32'd100173978);
    Send_IMC_Command(32'd93755920);
    Send_IMC_Command(32'd92868763);
    Send_IMC_Command(32'd93952792);
    Send_IMC_Command(32'd100374172);
    Send_IMC_Command(32'd92799133);
    Send_IMC_Command(32'd93953288);
    Send_IMC_Command(32'd93166750);
    Send_IMC_Command(32'd93232659);
    Send_IMC_Command(32'd95131551);
    Send_IMC_Command(32'd93298592);
    Send_IMC_Command(32'd93102083);
    Send_IMC_Command(32'd92459681);
    Send_IMC_Command(32'd93954466);
    Send_IMC_Command(32'd93429667);
    Send_IMC_Command(32'd93363364);
    Send_IMC_Command(32'd95062693);
    Send_IMC_Command(32'd93168898);
    Send_IMC_Command(32'd100305830);
    Send_IMC_Command(32'd93103634);
    Send_IMC_Command(32'd95025575);
    Send_IMC_Command(32'd94480304);
    Send_IMC_Command(32'd94810122);
    Send_IMC_Command(32'd94744602);
    Send_IMC_Command(32'd92379825);
    Send_IMC_Command(32'd100570034);
    Send_IMC_Command(32'd93630998);
    Send_IMC_Command(32'd95327667);
    Send_IMC_Command(32'd93500166);
    Send_IMC_Command(32'd92657076);
    Send_IMC_Command(32'd100571573);
    Send_IMC_Command(32'd97622198);
    Send_IMC_Command(32'd95260855);
    Send_IMC_Command(32'd93566725);
    Send_IMC_Command(32'd95204536);
    Send_IMC_Command(32'd100503993);
    Send_IMC_Command(32'd93501717);
    Send_IMC_Command(32'd100448442);
    Send_IMC_Command(32'd96057869);
    Send_IMC_Command(32'd95926813);
    Send_IMC_Command(32'd95392955);
    Send_IMC_Command(32'd93764359);
    Send_IMC_Command(32'd95335868);
    Send_IMC_Command(32'd96189471);
    Send_IMC_Command(32'd100636093);
    Send_IMC_Command(32'd96255247);
    Send_IMC_Command(32'd93830423);
    Send_IMC_Command(32'd93631678);
    Send_IMC_Command(32'd84327950);
    Send_IMC_Command(32'd94876095);
    Send_IMC_Command(32'd94093073);
    Send_IMC_Command(32'd93193152);
    Send_IMC_Command(32'd94552075);
    Send_IMC_Command(32'd92976833);
    Send_IMC_Command(32'd85508377);
    Send_IMC_Command(32'd93262786);
    Send_IMC_Command(32'd94552603);
    Send_IMC_Command(32'd97959619);
    Send_IMC_Command(32'd93569822);
    Send_IMC_Command(32'd97756356);
    Send_IMC_Command(32'd100451348);
    Send_IMC_Command(32'd92513221);
    Send_IMC_Command(32'd95208708);
    Send_IMC_Command(32'd93041094);
    Send_IMC_Command(32'd84461065);
    Send_IMC_Command(32'd94218183);
    Send_IMC_Command(32'd95864577);
    Send_IMC_Command(32'd92576200);
    Send_IMC_Command(32'd97765577);
    Send_IMC_Command(32'd94619916);
    Send_IMC_Command(32'd92513482);
    Send_IMC_Command(32'd93965003);
    Send_IMC_Command(32'd97831708);
    Send_IMC_Command(32'd83888264);
    Send_IMC_Command(32'd84940937);
    Send_IMC_Command(32'd83954058);
    Send_IMC_Command(32'd85006731);
    Send_IMC_Command(32'd84019852);
    Send_IMC_Command(32'd85072525);
    Send_IMC_Command(32'd84085646);
    Send_IMC_Command(32'd85138319);
    Send_IMC_Command(32'd84151440);
    Send_IMC_Command(32'd85204113);
    Send_IMC_Command(32'd84217234);
    Send_IMC_Command(32'd85269907);
    Send_IMC_Command(32'd84283028);
    Send_IMC_Command(32'd85335701);
    Send_IMC_Command(32'd85401494);
    Send_IMC_Command(32'd84348823);
    Send_IMC_Command(32'd84445592);
    Send_IMC_Command(32'd93821056);
    Send_IMC_Command(32'd84350873);
    Send_IMC_Command(32'd85493914);
    Send_IMC_Command(32'd93756112);
    Send_IMC_Command(32'd92917915);
    Send_IMC_Command(32'd93953016);
    Send_IMC_Command(32'd85694108);
    Send_IMC_Command(32'd92831901);
    Send_IMC_Command(32'd93953448);
    Send_IMC_Command(32'd93166750);
    Send_IMC_Command(32'd93232851);
    Send_IMC_Command(32'd84645791);
    Send_IMC_Command(32'd93298592);
    Send_IMC_Command(32'd93102211);
    Send_IMC_Command(32'd84021921);
    Send_IMC_Command(32'd93954466);
    Send_IMC_Command(32'd93429667);
    Send_IMC_Command(32'd93363364);
    Send_IMC_Command(32'd84576933);
    Send_IMC_Command(32'd93169026);
    Send_IMC_Command(32'd85625766);
    Send_IMC_Command(32'd93103826);
    Send_IMC_Command(32'd84482471);
    Send_IMC_Command(32'd94480304);
    Send_IMC_Command(32'd94810282);
    Send_IMC_Command(32'd94744826);
    Send_IMC_Command(32'd83991217);
    Send_IMC_Command(32'd85889970);
    Send_IMC_Command(32'd93631190);
    Send_IMC_Command(32'd84841907);
    Send_IMC_Command(32'd93500294);
    Send_IMC_Command(32'd84219316);
    Send_IMC_Command(32'd85891509);
    Send_IMC_Command(32'd85039286);
    Send_IMC_Command(32'd84775095);
    Send_IMC_Command(32'd93566853);
    Send_IMC_Command(32'd84718776);
    Send_IMC_Command(32'd85823929);
    Send_IMC_Command(32'd93501909);
    Send_IMC_Command(32'd85768378);
    Send_IMC_Command(32'd96058029);
    Send_IMC_Command(32'd95927037);
    Send_IMC_Command(32'd84907195);
    Send_IMC_Command(32'd93764487);
    Send_IMC_Command(32'd84850108);
    Send_IMC_Command(32'd96189695);
    Send_IMC_Command(32'd85956029);
    Send_IMC_Command(32'd96255407);
    Send_IMC_Command(32'd93830615);
    Send_IMC_Command(32'd93631678);
    Send_IMC_Command(32'd92716718);
    Send_IMC_Command(32'd94876095);
    Send_IMC_Command(32'd94093265);
    Send_IMC_Command(32'd93225920);
    Send_IMC_Command(32'd94552235);
    Send_IMC_Command(32'd92976833);
    Send_IMC_Command(32'd100188665);
    Send_IMC_Command(32'd93311938);
    Send_IMC_Command(32'd94552827);
    Send_IMC_Command(32'd85376707);
    Send_IMC_Command(32'd93570046);
    Send_IMC_Command(32'd85173444);
    Send_IMC_Command(32'd85771476);
    Send_IMC_Command(32'd84124613);
    Send_IMC_Command(32'd84723076);
    Send_IMC_Command(32'd93041094);
    Send_IMC_Command(32'd94946985);
    Send_IMC_Command(32'd94218183);
    Send_IMC_Command(32'd95864705);
    Send_IMC_Command(32'd84187592);
    Send_IMC_Command(32'd85182665);
    Send_IMC_Command(32'd94620076);
    Send_IMC_Command(32'd84124874);
    Send_IMC_Command(32'd93965003);
    Send_IMC_Command(32'd85249020);
    Send_IMC_Command(32'd85993608);
    Send_IMC_Command(32'd87046281);
    Send_IMC_Command(32'd86059402);
    Send_IMC_Command(32'd87112075);
    Send_IMC_Command(32'd86125196);
    Send_IMC_Command(32'd87177869);
    Send_IMC_Command(32'd86190990);
    Send_IMC_Command(32'd87243663);
    Send_IMC_Command(32'd86256784);
    Send_IMC_Command(32'd87309457);
    Send_IMC_Command(32'd86322578);
    Send_IMC_Command(32'd87375251);
    Send_IMC_Command(32'd86388372);
    Send_IMC_Command(32'd87441045);
    Send_IMC_Command(32'd87506838);
    Send_IMC_Command(32'd86454167);
    Send_IMC_Command(32'd86542768);
    Send_IMC_Command(32'd93827232);
    Send_IMC_Command(32'd86456241);
    Send_IMC_Command(32'd87591090);
    Send_IMC_Command(32'd93762288);
    Send_IMC_Command(32'd92926131);
    Send_IMC_Command(32'd95531928);
    Send_IMC_Command(32'd87791284);
    Send_IMC_Command(32'd92840117);
    Send_IMC_Command(32'd95532488);
    Send_IMC_Command(32'd93172918);
    Send_IMC_Command(32'd93239027);
    Send_IMC_Command(32'd86742967);
    Send_IMC_Command(32'd93304760);
    Send_IMC_Command(32'd93108387);
    Send_IMC_Command(32'd86127289);
    Send_IMC_Command(32'd95533498);
    Send_IMC_Command(32'd93435835);
    Send_IMC_Command(32'd93369532);
    Send_IMC_Command(32'd86674109);
    Send_IMC_Command(32'd93175202);
    Send_IMC_Command(32'd87722942);
    Send_IMC_Command(32'd93110002);
    Send_IMC_Command(32'd86587839);
    Send_IMC_Command(32'd96059328);
    Send_IMC_Command(32'd96387274);
    Send_IMC_Command(32'd96321690);
    Send_IMC_Command(32'd86094529);
    Send_IMC_Command(32'd87987138);
    Send_IMC_Command(32'd93635318);
    Send_IMC_Command(32'd86939075);
    Send_IMC_Command(32'd93504422);
    Send_IMC_Command(32'd86324676);
    Send_IMC_Command(32'd87994821);
    Send_IMC_Command(32'd87142598);
    Send_IMC_Command(32'd86872263);
    Send_IMC_Command(32'd93570981);
    Send_IMC_Command(32'd86820056);
    Send_IMC_Command(32'd87921113);
    Send_IMC_Command(32'd93510133);
    Send_IMC_Command(32'd87873754);
    Send_IMC_Command(32'd98163405);
    Send_IMC_Command(32'd96983709);
    Send_IMC_Command(32'd87004379);
    Send_IMC_Command(32'd93772711);
    Send_IMC_Command(32'd86951388);
    Send_IMC_Command(32'd98294943);
    Send_IMC_Command(32'd88053213);
    Send_IMC_Command(32'd98360783);
    Send_IMC_Command(32'd93838839);
    Send_IMC_Command(32'd93635806);
    Send_IMC_Command(32'd94822094);
    Send_IMC_Command(32'd96453087);
    Send_IMC_Command(32'd95674353);
    Send_IMC_Command(32'd93234144);
    Send_IMC_Command(32'd96133323);
    Send_IMC_Command(32'd92980961);
    Send_IMC_Command(32'd93905305);
    Send_IMC_Command(32'd93320162);
    Send_IMC_Command(32'd96133787);
    Send_IMC_Command(32'd87482083);
    Send_IMC_Command(32'd93578142);
    Send_IMC_Command(32'd87276772);
    Send_IMC_Command(32'd87876852);
    Send_IMC_Command(32'd86227941);
    Send_IMC_Command(32'd86828452);
    Send_IMC_Command(32'd93045222);
    Send_IMC_Command(32'd97052361);
    Send_IMC_Command(32'd95797223);
    Send_IMC_Command(32'd96921505);
    Send_IMC_Command(32'd86290920);
    Send_IMC_Command(32'd87288041);
    Send_IMC_Command(32'd96201164);
    Send_IMC_Command(32'd86228202);
    Send_IMC_Command(32'd95546091);
    Send_IMC_Command(32'd87354268);
    Send_IMC_Command(32'd94423176);
    Send_IMC_Command(32'd99653769);
    Send_IMC_Command(32'd94488970);
    Send_IMC_Command(32'd99719563);
    Send_IMC_Command(32'd94554764);
    Send_IMC_Command(32'd99785357);
    Send_IMC_Command(32'd94620558);
    Send_IMC_Command(32'd99851151);
    Send_IMC_Command(32'd94686352);
    Send_IMC_Command(32'd99916945);
    Send_IMC_Command(32'd94752146);
    Send_IMC_Command(32'd99982739);
    Send_IMC_Command(32'd94817940);
    Send_IMC_Command(32'd100048533);
    Send_IMC_Command(32'd100114326);
    Send_IMC_Command(32'd94883735);
    Send_IMC_Command(32'd97028528);
    Send_IMC_Command(32'd93827104);
    Send_IMC_Command(32'd94894001);
    Send_IMC_Command(32'd93882546);
    Send_IMC_Command(32'd93762096);
    Send_IMC_Command(32'd92876979);
    Send_IMC_Command(32'd95531832);
    Send_IMC_Command(32'd94082740);
    Send_IMC_Command(32'd92807349);
    Send_IMC_Command(32'd95532328);
    Send_IMC_Command(32'd93172918);
    Send_IMC_Command(32'd93238835);
    Send_IMC_Command(32'd97228727);
    Send_IMC_Command(32'd93304760);
    Send_IMC_Command(32'd93108259);
    Send_IMC_Command(32'd94565049);
    Send_IMC_Command(32'd95533498);
    Send_IMC_Command(32'd93435835);
    Send_IMC_Command(32'd93369532);
    Send_IMC_Command(32'd97159869);
    Send_IMC_Command(32'd93175074);
    Send_IMC_Command(32'd94014398);
    Send_IMC_Command(32'd93109810);
    Send_IMC_Command(32'd97098175);
    Send_IMC_Command(32'd96059328);
    Send_IMC_Command(32'd96387114);
    Send_IMC_Command(32'd96321594);
    Send_IMC_Command(32'd94483137);
    Send_IMC_Command(32'd94278594);
    Send_IMC_Command(32'd93635126);
    Send_IMC_Command(32'd97424835);
    Send_IMC_Command(32'd93504294);
    Send_IMC_Command(32'd94762436);
    Send_IMC_Command(32'd94286277);
    Send_IMC_Command(32'd99725510);
    Send_IMC_Command(32'd97358023);
    Send_IMC_Command(32'd93570853);
    Send_IMC_Command(32'd97305816);
    Send_IMC_Command(32'd94212569);
    Send_IMC_Command(32'd93509941);
    Send_IMC_Command(32'd94165210);
    Send_IMC_Command(32'd98163245);
    Send_IMC_Command(32'd96983613);
    Send_IMC_Command(32'd97490139);
    Send_IMC_Command(32'd93772583);
    Send_IMC_Command(32'd97437148);
    Send_IMC_Command(32'd98294847);
    Send_IMC_Command(32'd94344669);
    Send_IMC_Command(32'd98360623);
    Send_IMC_Command(32'd93838647);
    Send_IMC_Command(32'd93635806);
    Send_IMC_Command(32'd86433326);
    Send_IMC_Command(32'd96453087);
    Send_IMC_Command(32'd95674161);
    Send_IMC_Command(32'd93201376);
    Send_IMC_Command(32'd96133163);
    Send_IMC_Command(32'd92980961);
    Send_IMC_Command(32'd87613753);
    Send_IMC_Command(32'd93271010);
    Send_IMC_Command(32'd96133691);
    Send_IMC_Command(32'd100064995);
    Send_IMC_Command(32'd93578046);
    Send_IMC_Command(32'd99859684);
    Send_IMC_Command(32'd94168116);
    Send_IMC_Command(32'd94616549);
    Send_IMC_Command(32'd97314084);
    Send_IMC_Command(32'd93045222);
    Send_IMC_Command(32'd86566441);
    Send_IMC_Command(32'd95797223);
    Send_IMC_Command(32'd96921377);
    Send_IMC_Command(32'd94679528);
    Send_IMC_Command(32'd99870953);
    Send_IMC_Command(32'd96201004);
    Send_IMC_Command(32'd94616810);
    Send_IMC_Command(32'd95546091);
    Send_IMC_Command(32'd99937084);
    Send_IMC_Command(32'd85993608);
    Send_IMC_Command(32'd87046281);
    Send_IMC_Command(32'd86059402);
    Send_IMC_Command(32'd87112075);
    Send_IMC_Command(32'd86125196);
    Send_IMC_Command(32'd87177869);
    Send_IMC_Command(32'd86190990);
    Send_IMC_Command(32'd87243663);
    Send_IMC_Command(32'd86256784);
    Send_IMC_Command(32'd87309457);
    Send_IMC_Command(32'd86322578);
    Send_IMC_Command(32'd87375251);
    Send_IMC_Command(32'd86388372);
    Send_IMC_Command(32'd87441045);
    Send_IMC_Command(32'd87506838);
    Send_IMC_Command(32'd86454167);
    Send_IMC_Command(32'd86542768);
    Send_IMC_Command(32'd93827232);
    Send_IMC_Command(32'd86456241);
    Send_IMC_Command(32'd87591090);
    Send_IMC_Command(32'd93762288);
    Send_IMC_Command(32'd92926131);
    Send_IMC_Command(32'd95531928);
    Send_IMC_Command(32'd87791284);
    Send_IMC_Command(32'd92840117);
    Send_IMC_Command(32'd95532488);
    Send_IMC_Command(32'd93172918);
    Send_IMC_Command(32'd93239027);
    Send_IMC_Command(32'd86742967);
    Send_IMC_Command(32'd93304760);
    Send_IMC_Command(32'd93108387);
    Send_IMC_Command(32'd86127289);
    Send_IMC_Command(32'd95533498);
    Send_IMC_Command(32'd93435835);
    Send_IMC_Command(32'd93369532);
    Send_IMC_Command(32'd86674109);
    Send_IMC_Command(32'd93175202);
    Send_IMC_Command(32'd87722942);
    Send_IMC_Command(32'd93110002);
    Send_IMC_Command(32'd86587839);
    Send_IMC_Command(32'd96059328);
    Send_IMC_Command(32'd96387274);
    Send_IMC_Command(32'd96321690);
    Send_IMC_Command(32'd86094529);
    Send_IMC_Command(32'd87987138);
    Send_IMC_Command(32'd93635318);
    Send_IMC_Command(32'd86939075);
    Send_IMC_Command(32'd93504422);
    Send_IMC_Command(32'd86324676);
    Send_IMC_Command(32'd87994821);
    Send_IMC_Command(32'd87142598);
    Send_IMC_Command(32'd86872263);
    Send_IMC_Command(32'd93570981);
    Send_IMC_Command(32'd86820056);
    Send_IMC_Command(32'd87921113);
    Send_IMC_Command(32'd93510133);
    Send_IMC_Command(32'd87873754);
    Send_IMC_Command(32'd98163405);
    Send_IMC_Command(32'd96983709);
    Send_IMC_Command(32'd87004379);
    Send_IMC_Command(32'd93772711);
    Send_IMC_Command(32'd86951388);
    Send_IMC_Command(32'd98294943);
    Send_IMC_Command(32'd88053213);
    Send_IMC_Command(32'd98360783);
    Send_IMC_Command(32'd93838839);
    Send_IMC_Command(32'd93635806);
    Send_IMC_Command(32'd94822094);
    Send_IMC_Command(32'd96453087);
    Send_IMC_Command(32'd95674353);
    Send_IMC_Command(32'd93234144);
    Send_IMC_Command(32'd96133323);
    Send_IMC_Command(32'd92980961);
    Send_IMC_Command(32'd93905305);
    Send_IMC_Command(32'd93320162);
    Send_IMC_Command(32'd96133787);
    Send_IMC_Command(32'd87482083);
    Send_IMC_Command(32'd93578142);
    Send_IMC_Command(32'd87276772);
    Send_IMC_Command(32'd87876852);
    Send_IMC_Command(32'd86227941);
    Send_IMC_Command(32'd86828452);
    Send_IMC_Command(32'd93045222);
    Send_IMC_Command(32'd97052361);
    Send_IMC_Command(32'd95797223);
    Send_IMC_Command(32'd96921505);
    Send_IMC_Command(32'd86290920);
    Send_IMC_Command(32'd87288041);
    Send_IMC_Command(32'd96201164);
    Send_IMC_Command(32'd86228202);
    Send_IMC_Command(32'd95546091);
    Send_IMC_Command(32'd87354268);
    Send_IMC_Command(32'd88098952);
    Send_IMC_Command(32'd89151625);
    Send_IMC_Command(32'd88164746);
    Send_IMC_Command(32'd89217419);
    Send_IMC_Command(32'd88230540);
    Send_IMC_Command(32'd89283213);
    Send_IMC_Command(32'd88296334);
    Send_IMC_Command(32'd89349007);
    Send_IMC_Command(32'd88362160);
    Send_IMC_Command(32'd89414833);
    Send_IMC_Command(32'd88427954);
    Send_IMC_Command(32'd89480627);
    Send_IMC_Command(32'd88493748);
    Send_IMC_Command(32'd89546421);
    Send_IMC_Command(32'd89612214);
    Send_IMC_Command(32'd88559543);
    Send_IMC_Command(32'd88639960);
    Send_IMC_Command(32'd95934656);
    Send_IMC_Command(32'd88561625);
    Send_IMC_Command(32'd89688282);
    Send_IMC_Command(32'd95869584);
    Send_IMC_Command(32'd92901595);
    Send_IMC_Command(32'd98163640);
    Send_IMC_Command(32'd89896668);
    Send_IMC_Command(32'd92848349);
    Send_IMC_Command(32'd98164200);
    Send_IMC_Command(32'd93183198);
    Send_IMC_Command(32'd93249171);
    Send_IMC_Command(32'd88848351);
    Send_IMC_Command(32'd93315040);
    Send_IMC_Command(32'd93118659);
    Send_IMC_Command(32'd88232673);
    Send_IMC_Command(32'd98165218);
    Send_IMC_Command(32'd95543267);
    Send_IMC_Command(32'd95476964);
    Send_IMC_Command(32'd88771301);
    Send_IMC_Command(32'd93185474);
    Send_IMC_Command(32'd89820134);
    Send_IMC_Command(32'd93120146);
    Send_IMC_Command(32'd88693223);
    Send_IMC_Command(32'd98690816);
    Send_IMC_Command(32'd98959594);
    Send_IMC_Command(32'd98894010);
    Send_IMC_Command(32'd88201729);
    Send_IMC_Command(32'd90092290);
    Send_IMC_Command(32'd95683222);
    Send_IMC_Command(32'd89044227);
    Send_IMC_Command(32'd95552454);
    Send_IMC_Command(32'd88429828);
    Send_IMC_Command(32'd90102021);
    Send_IMC_Command(32'd89249798);
    Send_IMC_Command(32'd88977415);
    Send_IMC_Command(32'd95619013);
    Send_IMC_Command(32'd88867848);
    Send_IMC_Command(32'd90026249);
    Send_IMC_Command(32'd95553941);
    Send_IMC_Command(32'd89917450);
    Send_IMC_Command(32'd84478701);
    Send_IMC_Command(32'd84347581);
    Send_IMC_Command(32'd89109515);
    Send_IMC_Command(32'd95816647);
    Send_IMC_Command(32'd88999180);
    Send_IMC_Command(32'd84610239);
    Send_IMC_Command(32'd90158349);
    Send_IMC_Command(32'd84676079);
    Send_IMC_Command(32'd95882647);
    Send_IMC_Command(32'd95683598);
    Send_IMC_Command(32'd96866030);
    Send_IMC_Command(32'd99025167);
    Send_IMC_Command(32'd98242449);
    Send_IMC_Command(32'd93242128);
    Send_IMC_Command(32'd98701547);
    Send_IMC_Command(32'd92931601);
    Send_IMC_Command(32'd95949241);
    Send_IMC_Command(32'd93295378);
    Send_IMC_Command(32'd98702011);
    Send_IMC_Command(32'd89525779);
    Send_IMC_Command(32'd95622078);
    Send_IMC_Command(32'd89383956);
    Send_IMC_Command(32'd89920660);
    Send_IMC_Command(32'd88335125);
    Send_IMC_Command(32'd88872388);
    Send_IMC_Command(32'd92995862);
    Send_IMC_Command(32'd99096297);
    Send_IMC_Command(32'd98428695);
    Send_IMC_Command(32'd84285377);
    Send_IMC_Command(32'd88398104);
    Send_IMC_Command(32'd89331737);
    Send_IMC_Command(32'd98769388);
    Send_IMC_Command(32'd88335386);
    Send_IMC_Command(32'd98114075);
    Send_IMC_Command(32'd89398204);
    Send_IMC_Command(32'd96528520);
    Send_IMC_Command(32'd93370505);
    Send_IMC_Command(32'd96594314);
    Send_IMC_Command(32'd93436299);
    Send_IMC_Command(32'd96660108);
    Send_IMC_Command(32'd93502093);
    Send_IMC_Command(32'd96725902);
    Send_IMC_Command(32'd93567887);
    Send_IMC_Command(32'd96791728);
    Send_IMC_Command(32'd93633713);
    Send_IMC_Command(32'd96857522);
    Send_IMC_Command(32'd93699507);
    Send_IMC_Command(32'd96923316);
    Send_IMC_Command(32'd93765301);
    Send_IMC_Command(32'd93831094);
    Send_IMC_Command(32'd96989111);
    Send_IMC_Command(32'd99125720);
    Send_IMC_Command(32'd95934528);
    Send_IMC_Command(32'd96966617);
    Send_IMC_Command(32'd95979738);
    Send_IMC_Command(32'd95869520);
    Send_IMC_Command(32'd92885211);
    Send_IMC_Command(32'd98163544);
    Send_IMC_Command(32'd96188124);
    Send_IMC_Command(32'd92815581);
    Send_IMC_Command(32'd98164040);
    Send_IMC_Command(32'd93183198);
    Send_IMC_Command(32'd93249107);
    Send_IMC_Command(32'd99334111);
    Send_IMC_Command(32'd93315040);
    Send_IMC_Command(32'd93118531);
    Send_IMC_Command(32'd96637665);
    Send_IMC_Command(32'd98165218);
    Send_IMC_Command(32'd95543267);
    Send_IMC_Command(32'd95476964);
    Send_IMC_Command(32'd99257061);
    Send_IMC_Command(32'd93185346);
    Send_IMC_Command(32'd96111590);
    Send_IMC_Command(32'd93120082);
    Send_IMC_Command(32'd99203559);
    Send_IMC_Command(32'd98690816);
    Send_IMC_Command(32'd98959434);
    Send_IMC_Command(32'd98893914);
    Send_IMC_Command(32'd96590337);
    Send_IMC_Command(32'd96383746);
    Send_IMC_Command(32'd95683158);
    Send_IMC_Command(32'd99529987);
    Send_IMC_Command(32'd95552326);
    Send_IMC_Command(32'd96834820);
    Send_IMC_Command(32'd96393477);
    Send_IMC_Command(32'd93444102);
    Send_IMC_Command(32'd99463175);
    Send_IMC_Command(32'd95618885);
    Send_IMC_Command(32'd99353608);
    Send_IMC_Command(32'd96317705);
    Send_IMC_Command(32'd95553877);
    Send_IMC_Command(32'd96208906);
    Send_IMC_Command(32'd84478541);
    Send_IMC_Command(32'd84347485);
    Send_IMC_Command(32'd99595275);
    Send_IMC_Command(32'd95816519);
    Send_IMC_Command(32'd99484940);
    Send_IMC_Command(32'd84610143);
    Send_IMC_Command(32'd96449805);
    Send_IMC_Command(32'd84675919);
    Send_IMC_Command(32'd95882583);
    Send_IMC_Command(32'd95683598);
    Send_IMC_Command(32'd88477262);
    Send_IMC_Command(32'd99025167);
    Send_IMC_Command(32'd98242385);
    Send_IMC_Command(32'd93209360);
    Send_IMC_Command(32'd98701387);
    Send_IMC_Command(32'd92931601);
    Send_IMC_Command(32'd89657689);
    Send_IMC_Command(32'd93278994);
    Send_IMC_Command(32'd98701915);
    Send_IMC_Command(32'd93720083);
    Send_IMC_Command(32'd95621982);
    Send_IMC_Command(32'd93578260);
    Send_IMC_Command(32'd96212052);
    Send_IMC_Command(32'd96723733);
    Send_IMC_Command(32'd99358020);
    Send_IMC_Command(32'd92995862);
    Send_IMC_Command(32'd88610377);
    Send_IMC_Command(32'd98428695);
    Send_IMC_Command(32'd84285249);
    Send_IMC_Command(32'd96786712);
    Send_IMC_Command(32'd93526041);
    Send_IMC_Command(32'd98769228);
    Send_IMC_Command(32'd96723994);
    Send_IMC_Command(32'd98114075);
    Send_IMC_Command(32'd93592412);
    Send_IMC_Command(32'd88098952);
    Send_IMC_Command(32'd89151625);
    Send_IMC_Command(32'd88164746);
    Send_IMC_Command(32'd89217419);
    Send_IMC_Command(32'd88230540);
    Send_IMC_Command(32'd89283213);
    Send_IMC_Command(32'd88296334);
    Send_IMC_Command(32'd89349007);
    Send_IMC_Command(32'd88362160);
    Send_IMC_Command(32'd89414833);
    Send_IMC_Command(32'd88427954);
    Send_IMC_Command(32'd89480627);
    Send_IMC_Command(32'd88493748);
    Send_IMC_Command(32'd89546421);
    Send_IMC_Command(32'd89612214);
    Send_IMC_Command(32'd88559543);
    Send_IMC_Command(32'd88639960);
    Send_IMC_Command(32'd95934656);
    Send_IMC_Command(32'd88561625);
    Send_IMC_Command(32'd89688282);
    Send_IMC_Command(32'd95869584);
    Send_IMC_Command(32'd92901595);
    Send_IMC_Command(32'd98163640);
    Send_IMC_Command(32'd89896668);
    Send_IMC_Command(32'd92848349);
    Send_IMC_Command(32'd98164200);
    Send_IMC_Command(32'd93183198);
    Send_IMC_Command(32'd93249171);
    Send_IMC_Command(32'd88848351);
    Send_IMC_Command(32'd93315040);
    Send_IMC_Command(32'd93118659);
    Send_IMC_Command(32'd88232673);
    Send_IMC_Command(32'd98165218);
    Send_IMC_Command(32'd95543267);
    Send_IMC_Command(32'd95476964);
    Send_IMC_Command(32'd88771301);
    Send_IMC_Command(32'd93185474);
    Send_IMC_Command(32'd89820134);
    Send_IMC_Command(32'd93120146);
    Send_IMC_Command(32'd88693223);
    Send_IMC_Command(32'd98690816);
    Send_IMC_Command(32'd98959594);
    Send_IMC_Command(32'd98894010);
    Send_IMC_Command(32'd88201729);
    Send_IMC_Command(32'd90092290);
    Send_IMC_Command(32'd95683222);
    Send_IMC_Command(32'd89044227);
    Send_IMC_Command(32'd95552454);
    Send_IMC_Command(32'd88429828);
    Send_IMC_Command(32'd90102021);
    Send_IMC_Command(32'd89249798);
    Send_IMC_Command(32'd88977415);
    Send_IMC_Command(32'd95619013);
    Send_IMC_Command(32'd88867848);
    Send_IMC_Command(32'd90026249);
    Send_IMC_Command(32'd95553941);
    Send_IMC_Command(32'd89917450);
    Send_IMC_Command(32'd84478701);
    Send_IMC_Command(32'd84347581);
    Send_IMC_Command(32'd89109515);
    Send_IMC_Command(32'd95816647);
    Send_IMC_Command(32'd88999180);
    Send_IMC_Command(32'd84610239);
    Send_IMC_Command(32'd90158349);
    Send_IMC_Command(32'd84676079);
    Send_IMC_Command(32'd95882647);
    Send_IMC_Command(32'd95683598);
    Send_IMC_Command(32'd96866030);
    Send_IMC_Command(32'd99025167);
    Send_IMC_Command(32'd98242449);
    Send_IMC_Command(32'd93242128);
    Send_IMC_Command(32'd98701547);
    Send_IMC_Command(32'd92931601);
    Send_IMC_Command(32'd95949241);
    Send_IMC_Command(32'd93295378);
    Send_IMC_Command(32'd98702011);
    Send_IMC_Command(32'd89525779);
    Send_IMC_Command(32'd95622078);
    Send_IMC_Command(32'd89383956);
    Send_IMC_Command(32'd89920660);
    Send_IMC_Command(32'd88335125);
    Send_IMC_Command(32'd88872388);
    Send_IMC_Command(32'd92995862);
    Send_IMC_Command(32'd99096297);
    Send_IMC_Command(32'd98428695);
    Send_IMC_Command(32'd84285377);
    Send_IMC_Command(32'd88398104);
    Send_IMC_Command(32'd89331737);
    Send_IMC_Command(32'd98769388);
    Send_IMC_Command(32'd88335386);
    Send_IMC_Command(32'd98114075);
    Send_IMC_Command(32'd89398204);
    Send_IMC_Command(32'd90204160);
    Send_IMC_Command(32'd91256833);
    Send_IMC_Command(32'd90269954);
    Send_IMC_Command(32'd91322627);
    Send_IMC_Command(32'd90335748);
    Send_IMC_Command(32'd91388421);
    Send_IMC_Command(32'd90401542);
    Send_IMC_Command(32'd91454215);
    Send_IMC_Command(32'd90467336);
    Send_IMC_Command(32'd91520009);
    Send_IMC_Command(32'd90533130);
    Send_IMC_Command(32'd91585803);
    Send_IMC_Command(32'd90598924);
    Send_IMC_Command(32'd91651597);
    Send_IMC_Command(32'd91717390);
    Send_IMC_Command(32'd90664719);
    Send_IMC_Command(32'd90702096);
    Send_IMC_Command(32'd84873440);
    Send_IMC_Command(32'd90666769);
    Send_IMC_Command(32'd91750418);
    Send_IMC_Command(32'd84808368);
    Send_IMC_Command(32'd83996691);
    Send_IMC_Command(32'd85005272);
    Send_IMC_Command(32'd91950612);
    Send_IMC_Command(32'd83943445);
    Send_IMC_Command(32'd85005704);
    Send_IMC_Command(32'd84218902);
    Send_IMC_Command(32'd84285107);
    Send_IMC_Command(32'd90902295);
    Send_IMC_Command(32'd84350744);
    Send_IMC_Command(32'd84154595);
    Send_IMC_Command(32'd90337817);
    Send_IMC_Command(32'd85006618);
    Send_IMC_Command(32'd84481819);
    Send_IMC_Command(32'd84415516);
    Send_IMC_Command(32'd90833437);
    Send_IMC_Command(32'd84221410);
    Send_IMC_Command(32'd91882270);
    Send_IMC_Command(32'd84156082);
    Send_IMC_Command(32'd90798367);
    Send_IMC_Command(32'd85532448);
    Send_IMC_Command(32'd85860490);
    Send_IMC_Command(32'd85795034);
    Send_IMC_Command(32'd90247713);
    Send_IMC_Command(32'd92146466);
    Send_IMC_Command(32'd84681398);
    Send_IMC_Command(32'd91098403);
    Send_IMC_Command(32'd84550630);
    Send_IMC_Command(32'd90535204);
    Send_IMC_Command(32'd92148005);
    Send_IMC_Command(32'd91295782);
    Send_IMC_Command(32'd91031591);
    Send_IMC_Command(32'd84617189);
    Send_IMC_Command(32'd90973224);
    Send_IMC_Command(32'd92080425);
    Send_IMC_Command(32'd84552117);
    Send_IMC_Command(32'd92022826);
    Send_IMC_Command(32'd86583949);
    Send_IMC_Command(32'd86452957);
    Send_IMC_Command(32'd91163691);
    Send_IMC_Command(32'd84814823);
    Send_IMC_Command(32'd91104556);
    Send_IMC_Command(32'd86715615);
    Send_IMC_Command(32'd92212525);
    Send_IMC_Command(32'd86781327);
    Send_IMC_Command(32'd84880823);
    Send_IMC_Command(32'd84681774);
    Send_IMC_Command(32'd98971278);
    Send_IMC_Command(32'd85926191);
    Send_IMC_Command(32'd85143473);
    Send_IMC_Command(32'd84337456);
    Send_IMC_Command(32'd85602443);
    Send_IMC_Command(32'd84026929);
    Send_IMC_Command(32'd98054617);
    Send_IMC_Command(32'd84390706);
    Send_IMC_Command(32'd85603035);
    Send_IMC_Command(32'd91631155);
    Send_IMC_Command(32'd84620254);
    Send_IMC_Command(32'd91429940);
    Send_IMC_Command(32'd92026036);
    Send_IMC_Command(32'd90381109);
    Send_IMC_Command(32'd90977764);
    Send_IMC_Command(32'd84091190);
    Send_IMC_Command(32'd92812937);
    Send_IMC_Command(32'd85270327);
    Send_IMC_Command(32'd86390753);
    Send_IMC_Command(32'd90444088);
    Send_IMC_Command(32'd91437113);
    Send_IMC_Command(32'd85670284);
    Send_IMC_Command(32'd90381370);
    Send_IMC_Command(32'd85015099);
    Send_IMC_Command(32'd91503580);
    Send_IMC_Command(32'd98600960);
    Send_IMC_Command(32'd95475713);
    Send_IMC_Command(32'd98666754);
    Send_IMC_Command(32'd95541507);
    Send_IMC_Command(32'd98732548);
    Send_IMC_Command(32'd95607301);
    Send_IMC_Command(32'd98798342);
    Send_IMC_Command(32'd95673095);
    Send_IMC_Command(32'd98864136);
    Send_IMC_Command(32'd95738889);
    Send_IMC_Command(32'd98929930);
    Send_IMC_Command(32'd95804683);
    Send_IMC_Command(32'd98995724);
    Send_IMC_Command(32'd95870477);
    Send_IMC_Command(32'd95936270);
    Send_IMC_Command(32'd99061519);
    Send_IMC_Command(32'd92799248);
    Send_IMC_Command(32'd84873312);
    Send_IMC_Command(32'd99071761);
    Send_IMC_Command(32'd98041874);
    Send_IMC_Command(32'd84808304);
    Send_IMC_Command(32'd83980307);
    Send_IMC_Command(32'd85005176);
    Send_IMC_Command(32'd98242068);
    Send_IMC_Command(32'd83910677);
    Send_IMC_Command(32'd85005672);
    Send_IMC_Command(32'd84218902);
    Send_IMC_Command(32'd84285043);
    Send_IMC_Command(32'd92999447);
    Send_IMC_Command(32'd84350744);
    Send_IMC_Command(32'd84154467);
    Send_IMC_Command(32'd98742809);
    Send_IMC_Command(32'd85006618);
    Send_IMC_Command(32'd84481819);
    Send_IMC_Command(32'd84415516);
    Send_IMC_Command(32'd92930589);
    Send_IMC_Command(32'd84221282);
    Send_IMC_Command(32'd98173726);
    Send_IMC_Command(32'd84156018);
    Send_IMC_Command(32'd92920095);
    Send_IMC_Command(32'd85532448);
    Send_IMC_Command(32'd85860458);
    Send_IMC_Command(32'd85794938);
    Send_IMC_Command(32'd98636321);
    Send_IMC_Command(32'd98437922);
    Send_IMC_Command(32'd84681334);
    Send_IMC_Command(32'd93195555);
    Send_IMC_Command(32'd84550502);
    Send_IMC_Command(32'd98940196);
    Send_IMC_Command(32'd98439461);
    Send_IMC_Command(32'd95490086);
    Send_IMC_Command(32'd93128743);
    Send_IMC_Command(32'd84617061);
    Send_IMC_Command(32'd93070376);
    Send_IMC_Command(32'd98371881);
    Send_IMC_Command(32'd84552053);
    Send_IMC_Command(32'd98314282);
    Send_IMC_Command(32'd86583917);
    Send_IMC_Command(32'd86452861);
    Send_IMC_Command(32'd93260843);
    Send_IMC_Command(32'd84814695);
    Send_IMC_Command(32'd93201708);
    Send_IMC_Command(32'd86715519);
    Send_IMC_Command(32'd98503981);
    Send_IMC_Command(32'd86781295);
    Send_IMC_Command(32'd84880759);
    Send_IMC_Command(32'd84681774);
    Send_IMC_Command(32'd90582638);
    Send_IMC_Command(32'd85926191);
    Send_IMC_Command(32'd85143409);
    Send_IMC_Command(32'd84304688);
    Send_IMC_Command(32'd85602411);
    Send_IMC_Command(32'd84026929);
    Send_IMC_Command(32'd91763065);
    Send_IMC_Command(32'd84374322);
    Send_IMC_Command(32'd85602939);
    Send_IMC_Command(32'd95825459);
    Send_IMC_Command(32'd84620158);
    Send_IMC_Command(32'd95624244);
    Send_IMC_Command(32'd98317428);
    Send_IMC_Command(32'd98769717);
    Send_IMC_Command(32'd93074788);
    Send_IMC_Command(32'd84091190);
    Send_IMC_Command(32'd90715753);
    Send_IMC_Command(32'd85270327);
    Send_IMC_Command(32'd86390625);
    Send_IMC_Command(32'd98832696);
    Send_IMC_Command(32'd95631417);
    Send_IMC_Command(32'd85670252);
    Send_IMC_Command(32'd98769978);
    Send_IMC_Command(32'd85015099);
    Send_IMC_Command(32'd95697788);
    Send_IMC_Command(32'd90204160);
    Send_IMC_Command(32'd91256833);
    Send_IMC_Command(32'd90269954);
    Send_IMC_Command(32'd91322627);
    Send_IMC_Command(32'd90335748);
    Send_IMC_Command(32'd91388421);
    Send_IMC_Command(32'd90401542);
    Send_IMC_Command(32'd91454215);
    Send_IMC_Command(32'd90467336);
    Send_IMC_Command(32'd91520009);
    Send_IMC_Command(32'd90533130);
    Send_IMC_Command(32'd91585803);
    Send_IMC_Command(32'd90598924);
    Send_IMC_Command(32'd91651597);
    Send_IMC_Command(32'd91717390);
    Send_IMC_Command(32'd90664719);
    Send_IMC_Command(32'd90702096);
    Send_IMC_Command(32'd84873440);
    Send_IMC_Command(32'd90666769);
    Send_IMC_Command(32'd91750418);
    Send_IMC_Command(32'd84808368);
    Send_IMC_Command(32'd83996691);
    Send_IMC_Command(32'd85005272);
    Send_IMC_Command(32'd91950612);
    Send_IMC_Command(32'd83943445);
    Send_IMC_Command(32'd85005704);
    Send_IMC_Command(32'd84218902);
    Send_IMC_Command(32'd84285107);
    Send_IMC_Command(32'd90902295);
    Send_IMC_Command(32'd84350744);
    Send_IMC_Command(32'd84154595);
    Send_IMC_Command(32'd90337817);
    Send_IMC_Command(32'd85006618);
    Send_IMC_Command(32'd84481819);
    Send_IMC_Command(32'd84415516);
    Send_IMC_Command(32'd90833437);
    Send_IMC_Command(32'd84221410);
    Send_IMC_Command(32'd91882270);
    Send_IMC_Command(32'd84156082);
    Send_IMC_Command(32'd90798367);
    Send_IMC_Command(32'd85532448);
    Send_IMC_Command(32'd85860490);
    Send_IMC_Command(32'd85795034);
    Send_IMC_Command(32'd90247713);
    Send_IMC_Command(32'd92146466);
    Send_IMC_Command(32'd84681398);
    Send_IMC_Command(32'd91098403);
    Send_IMC_Command(32'd84550630);
    Send_IMC_Command(32'd90535204);
    Send_IMC_Command(32'd92148005);
    Send_IMC_Command(32'd91295782);
    Send_IMC_Command(32'd91031591);
    Send_IMC_Command(32'd84617189);
    Send_IMC_Command(32'd90973224);
    Send_IMC_Command(32'd92080425);
    Send_IMC_Command(32'd84552117);
    Send_IMC_Command(32'd92022826);
    Send_IMC_Command(32'd86583949);
    Send_IMC_Command(32'd86452957);
    Send_IMC_Command(32'd91163691);
    Send_IMC_Command(32'd84814823);
    Send_IMC_Command(32'd91104556);
    Send_IMC_Command(32'd86715615);
    Send_IMC_Command(32'd92212525);
    Send_IMC_Command(32'd86781327);
    Send_IMC_Command(32'd84880823);
    Send_IMC_Command(32'd84681774);
    Send_IMC_Command(32'd98971278);
    Send_IMC_Command(32'd85926191);
    Send_IMC_Command(32'd85143473);
    Send_IMC_Command(32'd84337456);
    Send_IMC_Command(32'd85602443);
    Send_IMC_Command(32'd84026929);
    Send_IMC_Command(32'd98054617);
    Send_IMC_Command(32'd84390706);
    Send_IMC_Command(32'd85603035);
    Send_IMC_Command(32'd91631155);
    Send_IMC_Command(32'd84620254);
    Send_IMC_Command(32'd91429940);
    Send_IMC_Command(32'd92026036);
    Send_IMC_Command(32'd90381109);
    Send_IMC_Command(32'd90977764);
    Send_IMC_Command(32'd84091190);
    Send_IMC_Command(32'd92812937);
    Send_IMC_Command(32'd85270327);
    Send_IMC_Command(32'd86390753);
    Send_IMC_Command(32'd90444088);
    Send_IMC_Command(32'd91437113);
    Send_IMC_Command(32'd85670284);
    Send_IMC_Command(32'd90381370);
    Send_IMC_Command(32'd85015099);
    Send_IMC_Command(32'd91503580);

endtask