`timescale 1ns/1ps

module BCIM_tb;

import avalon_mm_pkg::*;
import verbosity_pkg::*;

import BCIM_PKG::*;


logic clk;
logic rst;

logic [7:0] stimulus;

logic [31:0] avalon_mm_addr;

logic [31:0] avalon_mm_wdata;
logic [31:0] avalon_mm_rdata;

logic       avalon_mm_waitreq, avalon_mm_readdatavalid, avalon_mm_read, avalon_mm_write;

logic [31:0] rd;

logic [7:0] state_bytes [15:0];
logic [7:0] plain_text_bytes [15:0];
logic [7:0] round_key_bytes [15:0];
logic [7:0] key_bytes [9:0][15:0];


localparam PIM_ADDR_BITS = 8;
localparam LOAD_OFFSET = 2**PIM_ADDR_BITS;

avalon_mm_sim_block avalon_mm_sim_block_inst (
    .clk               (clk), // clk.clk
    .reset             (rst), // clk_reset.reset
    .avm_address       (avalon_mm_addr), // m0.address
    .avm_readdata      (avalon_mm_rdata), // .readdata
    .avm_writedata     (avalon_mm_wdata), // .writedata
    .avm_waitrequest   (avalon_mm_waitreq), // .waitrequest
    .avm_write         (avalon_mm_write), // .write
    .avm_read          (avalon_mm_read), // .read
    .avm_readdatavalid (avalon_mm_readdatavalid) // .readdatavalid
);



prime_datapath prime_datapath_inst (
    .sys_clk_in                 (clk),
    .sys_reset_in               (rst),

    //IMC Main Master
    .IMC_mm_waitrequest_out     (avalon_mm_waitreq),
    .IMC_mm_readdata_out        (avalon_mm_rdata),
    .IMC_mm_readdatavalid_out   (avalon_mm_readdatavalid),

    .IMC_mm_writedata_in        (avalon_mm_wdata),
    .IMC_mm_address_in          (avalon_mm_addr[8:0]),
    .IMC_mm_write_in            (avalon_mm_write),
    .IMC_mm_read_in             (avalon_mm_read)
);



class tb_BCIM_class #(
    int ARRAY_WIDTH = 8, 
    int BUS_DATA_WIDTH
) extends BCIM_class#(
    .ARRAY_WIDTH(ARRAY_WIDTH),
    .BUS_DATA_WIDTH(BUS_DATA_WIDTH)
);

    function new(input string my_name, input string prgm);
        super.new(my_name, prgm);
    endfunction
    
    //"Harness" connecting virtual function from parent to TB implementation details
    function get_memory_array(input int addr, output [ARRAY_WIDTH-1:0] data);
        data = prime_datapath_inst.ram_model_inst.mem[addr];
    endfunction
    
    //"Harness" connecting virtual function from parent to TB implementation details
    // This task operates the bfm to read IMC data
    task read_memory_array(input int read_addr, output [ARRAY_WIDTH-1:0] rdata);
    
        avalon_mm_sim_block_inst.mm_master_bfm_0.set_command_address(read_addr);
        avalon_mm_sim_block_inst.mm_master_bfm_0.set_command_request(REQ_READ);
        
        avalon_mm_sim_block_inst.mm_master_bfm_0.push_command();
    
        @(negedge(avalon_mm_readdatavalid));
        
        avalon_mm_sim_block_inst.mm_master_bfm_0.pop_response();
        rdata = avalon_mm_sim_block_inst.mm_master_bfm_0.get_response_data(0);
    
    endtask
    
    //"Harness" connecting virtual function from parent to TB implementation details
    // This task operates the bfm to send IMC commands
    task send_imc_command(input [BUS_DATA_WIDTH-1:0] write_data);

        avalon_mm_sim_block_inst.mm_master_bfm_0.set_command_data(write_data,0); // Set index to zero for now
        avalon_mm_sim_block_inst.mm_master_bfm_0.set_command_address(0);
        avalon_mm_sim_block_inst.mm_master_bfm_0.set_command_request(REQ_WRITE);
    
        avalon_mm_sim_block_inst.mm_master_bfm_0.push_command();
        
        @(negedge(avalon_mm_write));
        avalon_mm_sim_block_inst.mm_master_bfm_0.pop_response();
        
        wait(prime_datapath_inst.rw_control_inst.state == 8'h1F);
        
    endtask

endclass


BCIM_class#(32,32) cipher_obj;
tb_BCIM_class#(32,32) tb_cipher_obj;

initial begin
    rst = 1'b1;
    $display("-- Simulation Starting (%t)ps --",$time);
    
    //verbosity_pkg::set_verbosity(VERBOSITY_DEBUG);
    
    #1us;
    rst = 1'b0;
    #1us;
    
    
    //set_command
    
    //Init BFM
    $display("Version %S",avalon_mm_sim_block_inst.mm_master_bfm_0.get_version());
    avalon_mm_sim_block_inst.mm_master_bfm_0.init();


    Compact_AES();
    inv_Compact_AES();
    
    cipher_obj = new("ECB_AES_parent", "ECB_AES");
    tb_cipher_obj = new("ECB_AES_child", "ECB_AES");
    
    cipher_obj.test_case_access(1);
    tb_cipher_obj.test_case_access(1);
    
    cipher_obj.test_write_sequence();
    tb_cipher_obj.test_write_sequence();
    
    //cipher_obj.read_memory_array(1,rd);
    //$display("%h",rd);
    //tb_cipher_obj.read_memory_array(1,rd);
    //$display("%h",rd);
    //tb_cipher_obj.get_memory_array(1,rd);
    //$display("%h",rd);
    
    cipher_obj.run_cipher();
    tb_cipher_obj.run_cipher();
    

    #128000;

    $display("-- Simulation Completed (%t)ps --",$time);
    $stop;
    #100;
end


initial begin
    clk = 1'b0;
    forever #42 clk = ~clk;

end

//-----------------------------------------------------------------------------------------------------------------
//                                              Tasks
//-----------------------------------------------------------------------------------------------------------------

task Avalon_MM_Bus_Write(input logic [31:0] write_addr, input logic [31:0] write_data);
    begin
        //$display("-- Sending Write Command (%t)ps --",$time);
        avalon_mm_sim_block_inst.mm_master_bfm_0.set_command_data(write_data,0); // Set index to zero for now
        avalon_mm_sim_block_inst.mm_master_bfm_0.set_command_address(write_addr);
        avalon_mm_sim_block_inst.mm_master_bfm_0.set_command_request(REQ_WRITE);
    
        avalon_mm_sim_block_inst.mm_master_bfm_0.push_command();
        
        @(negedge(avalon_mm_write));
        avalon_mm_sim_block_inst.mm_master_bfm_0.pop_response();
        
        //#1000ns;
    end
endtask

task PIM_Command(input logic [31:0] write_data);
    begin
        //$display("-- Sending Write Command (%t)ps --",$time);
        avalon_mm_sim_block_inst.mm_master_bfm_0.set_command_data(write_data,0); // Set index to zero for now
        avalon_mm_sim_block_inst.mm_master_bfm_0.set_command_address(0);
        avalon_mm_sim_block_inst.mm_master_bfm_0.set_command_request(REQ_WRITE);
    
        avalon_mm_sim_block_inst.mm_master_bfm_0.push_command();
        
        @(negedge(avalon_mm_write));
        avalon_mm_sim_block_inst.mm_master_bfm_0.pop_response();
        
        wait(prime_datapath_inst.rw_control_inst.state == 8'h1F);
        //#1000ns;
    end
endtask

task Avalon_MM_Bus_Read(input logic [31:0] read_addr, output logic [31:0] read_data);
    begin
    avalon_mm_sim_block_inst.mm_master_bfm_0.set_command_address(read_addr);
    avalon_mm_sim_block_inst.mm_master_bfm_0.set_command_request(REQ_READ);
    
    avalon_mm_sim_block_inst.mm_master_bfm_0.push_command();

    @(negedge(avalon_mm_readdatavalid));
    
    avalon_mm_sim_block_inst.mm_master_bfm_0.pop_response();
    read_data = avalon_mm_sim_block_inst.mm_master_bfm_0.get_response_data(0);
    end
endtask

task Load_Byte_PIM(input logic [7:0] byte_in, input logic [31:0] start_addr);

    @(posedge(clk));
    @(posedge(clk));
    $display("-- Loading %2h on WL %3h - %3h (%t)ps --",byte_in,start_addr,start_addr+7,$time);
    
    begin
        for (int i = 0; i < 8; i++) begin
            Avalon_MM_Bus_Write(start_addr+i+LOAD_OFFSET,byte_in[i]);
        end
    end
endtask


task Load_State_Bytes_1Col(input logic [7:0] byte_in [15:0], input logic [31:0] start_addr);
    Load_Byte_PIM(byte_in[15],start_addr+'h0);
    Load_Byte_PIM(byte_in[11],start_addr+'h8);
    Load_Byte_PIM(byte_in[7],start_addr+'h10);
    Load_Byte_PIM(byte_in[3],start_addr+'h18);

    Load_Byte_PIM(byte_in[14],start_addr+'h20);
    Load_Byte_PIM(byte_in[10],start_addr+'h28);
    Load_Byte_PIM(byte_in[6],start_addr+'h30);
    Load_Byte_PIM(byte_in[2],start_addr+'h38);

    Load_Byte_PIM(byte_in[13],start_addr+'h40);
    Load_Byte_PIM(byte_in[9],start_addr+'h48);
    Load_Byte_PIM(byte_in[5],start_addr+'h50);
    Load_Byte_PIM(byte_in[1],start_addr+'h58);

    Load_Byte_PIM(byte_in[12],start_addr+'h60);
    Load_Byte_PIM(byte_in[8],start_addr+'h68);
    Load_Byte_PIM(byte_in[4],start_addr+'h70);
    Load_Byte_PIM(byte_in[0],start_addr+'h78);
endtask





task Print_State_Bytes_1Col(input logic [31:0] start_addr, string tag);
    logic [7:0] state_bytes [15:0];
    
    wait(prime_datapath_inst.rw_control_inst.state == 8'h1F);
    @(posedge(clk));
    @(posedge(clk));
    
    
    for (int j = 0; j < 16; j++) begin
        for (int i = 0; i < 8; i++) begin
            state_bytes[j][i] = prime_datapath_inst.ram_model_inst.mem[start_addr+(j*8)+i][0];
        end
    end
    $display("---------------------");
    $display("\t%S",tag);
    $display("---------------------");
    $display("| %H | %H | %H | %H |",state_bytes[0],state_bytes[4],state_bytes[8],state_bytes[12]);
    $display("---------------------");
    $display("| %H | %H | %H | %H |",state_bytes[1],state_bytes[5],state_bytes[9],state_bytes[13]);
    $display("---------------------");
    $display("| %H | %H | %H | %H |",state_bytes[2],state_bytes[6],state_bytes[10],state_bytes[14]);
    $display("---------------------");
    $display("| %H | %H | %H | %H |",state_bytes[3],state_bytes[7],state_bytes[11],state_bytes[15]);
    $display("---------------------");
    
endtask



//-----------------------------------------------------------------------------------------------------------------
//                                              Intrinsics
//-----------------------------------------------------------------------------------------------------------------

task Compact_AES();
    //Load Plain Text
    //Column-Wise 0-3
    plain_text_bytes    = '{8'h32,8'h88,8'h31,8'hE0,  //Row 0
                            8'h43,8'h5A,8'h31,8'h37,
                            8'hF6,8'h30,8'h98,8'h07,
                            8'hA8,8'h8D,8'hA2,8'h34}; //Row 3
    Load_State_Bytes_1Col(plain_text_bytes,'h0);
    
    //#10us;
    //Print_State_Bytes_1Col('h0,"Plain Text:");
    
    
    round_key_bytes = '{8'h2B,8'h28,8'hAB,8'h09,  //Row 0
                        8'h7E,8'hAE,8'hF7,8'hCF,
                        8'h15,8'hD2,8'h15,8'h4F,
                        8'h16,8'hA6,8'h88,8'h3C}; //Row 3
    Load_State_Bytes_1Col(round_key_bytes,'h80);
    
    //#10us;
    //Print_State_Bytes_1Col('h80,"Initial Key");
    
    ARK();
    
    //#10us;
    //Print_State_Bytes_1Col('h00,"Initial Add Key");
    
    
    
    SBOX();
    
    //#10us;
    //Print_State_Bytes_1Col('h00,"Initial Add Key");
    
    MC();
    
    //#10us;
    //Print_State_Bytes_1Col('h80,"1 Col");
    
    
    
    key_bytes[0] = '{8'hA0,8'h88,8'h23,8'h2A,  //Row 0
                    8'hFA,8'h54,8'hA3,8'h6C,
                    8'hFE,8'h2C,8'h39,8'h76,
                    8'h17,8'hB1,8'h39,8'h05}; //Row 3
    Load_State_Bytes_1Col(key_bytes[0],'h00);
    
    
    ARK();
    
    #10us;
    Print_State_Bytes_1Col('h00,"Add Key 1");

endtask



task inv_Compact_AES();

    key_bytes[0] = '{8'hA0,8'h88,8'h23,8'h2A,  //Row 0
                    8'hFA,8'h54,8'hA3,8'h6C,
                    8'hFE,8'h2C,8'h39,8'h76,
                    8'h17,8'hB1,8'h39,8'h05}; //Row 3
    Load_State_Bytes_1Col(key_bytes[0],'h80);
    
    
    ARK();
    
    #10us;
    Print_State_Bytes_1Col('h00,"Inv Add Key 1");
    
    
    inv_MC();
    
    #10us;
    Print_State_Bytes_1Col('h80,"Inv Mix Cols");
    
    
    inv_SBOX();
    
    #10us;
    Print_State_Bytes_1Col('h80,"Inv SBOX");
    
    round_key_bytes = '{8'h2B,8'h28,8'hAB,8'h09,  //Row 0
                        8'h7E,8'hAE,8'hF7,8'hCF,
                        8'h15,8'hD2,8'h15,8'h4F,
                        8'h16,8'hA6,8'h88,8'h3C}; //Row 3
    Load_State_Bytes_1Col(round_key_bytes,'h00);
    
    
    ARK();
    
    #10us;
    Print_State_Bytes_1Col('h00,"Plaintext");


endtask




task ARK();
//State Input   00-7F
//Key Input     80-FF
//Output        00-7F

PIM_Command(32'd83918848);
PIM_Command(32'd83984641);
PIM_Command(32'd84050434);
PIM_Command(32'd84116227);
PIM_Command(32'd84182020);
PIM_Command(32'd84247813);
PIM_Command(32'd84313606);
PIM_Command(32'd84379399);
PIM_Command(32'd84445192);
PIM_Command(32'd84510985);
PIM_Command(32'd84576778);
PIM_Command(32'd84642571);
PIM_Command(32'd84708364);
PIM_Command(32'd84774157);
PIM_Command(32'd84839950);
PIM_Command(32'd84905743);
PIM_Command(32'd84971536);
PIM_Command(32'd85037329);
PIM_Command(32'd85103122);
PIM_Command(32'd85168915);
PIM_Command(32'd85234708);
PIM_Command(32'd85300501);
PIM_Command(32'd85366294);
PIM_Command(32'd85432087);
PIM_Command(32'd85497880);
PIM_Command(32'd85563673);
PIM_Command(32'd85629466);
PIM_Command(32'd85695259);
PIM_Command(32'd85761052);
PIM_Command(32'd85826845);
PIM_Command(32'd85892638);
PIM_Command(32'd85958431);
PIM_Command(32'd86024224);
PIM_Command(32'd86090017);
PIM_Command(32'd86155810);
PIM_Command(32'd86221603);
PIM_Command(32'd86287396);
PIM_Command(32'd86353189);
PIM_Command(32'd86418982);
PIM_Command(32'd86484775);
PIM_Command(32'd86550568);
PIM_Command(32'd86616361);
PIM_Command(32'd86682154);
PIM_Command(32'd86747947);
PIM_Command(32'd86813740);
PIM_Command(32'd86879533);
PIM_Command(32'd86945326);
PIM_Command(32'd87011119);
PIM_Command(32'd87076912);
PIM_Command(32'd87142705);
PIM_Command(32'd87208498);
PIM_Command(32'd87274291);
PIM_Command(32'd87340084);
PIM_Command(32'd87405877);
PIM_Command(32'd87471670);
PIM_Command(32'd87537463);
PIM_Command(32'd87603256);
PIM_Command(32'd87669049);
PIM_Command(32'd87734842);
PIM_Command(32'd87800635);
PIM_Command(32'd87866428);
PIM_Command(32'd87932221);
PIM_Command(32'd87998014);
PIM_Command(32'd88063807);
PIM_Command(32'd88129600);
PIM_Command(32'd88195393);
PIM_Command(32'd88261186);
PIM_Command(32'd88326979);
PIM_Command(32'd88392772);
PIM_Command(32'd88458565);
PIM_Command(32'd88524358);
PIM_Command(32'd88590151);
PIM_Command(32'd88655944);
PIM_Command(32'd88721737);
PIM_Command(32'd88787530);
PIM_Command(32'd88853323);
PIM_Command(32'd88919116);
PIM_Command(32'd88984909);
PIM_Command(32'd89050702);
PIM_Command(32'd89116495);
PIM_Command(32'd89182288);
PIM_Command(32'd89248081);
PIM_Command(32'd89313874);
PIM_Command(32'd89379667);
PIM_Command(32'd89445460);
PIM_Command(32'd89511253);
PIM_Command(32'd89577046);
PIM_Command(32'd89642839);
PIM_Command(32'd89708632);
PIM_Command(32'd89774425);
PIM_Command(32'd89840218);
PIM_Command(32'd89906011);
PIM_Command(32'd89971804);
PIM_Command(32'd90037597);
PIM_Command(32'd90103390);
PIM_Command(32'd90169183);
PIM_Command(32'd90234976);
PIM_Command(32'd90300769);
PIM_Command(32'd90366562);
PIM_Command(32'd90432355);
PIM_Command(32'd90498148);
PIM_Command(32'd90563941);
PIM_Command(32'd90629734);
PIM_Command(32'd90695527);
PIM_Command(32'd90761320);
PIM_Command(32'd90827113);
PIM_Command(32'd90892906);
PIM_Command(32'd90958699);
PIM_Command(32'd91024492);
PIM_Command(32'd91090285);
PIM_Command(32'd91156078);
PIM_Command(32'd91221871);
PIM_Command(32'd91287664);
PIM_Command(32'd91353457);
PIM_Command(32'd91419250);
PIM_Command(32'd91485043);
PIM_Command(32'd91550836);
PIM_Command(32'd91616629);
PIM_Command(32'd91682422);
PIM_Command(32'd91748215);
PIM_Command(32'd91814008);
PIM_Command(32'd91879801);
PIM_Command(32'd91945594);
PIM_Command(32'd92011387);
PIM_Command(32'd92077180);
PIM_Command(32'd92142973);
PIM_Command(32'd92208766);
PIM_Command(32'd92274559);


endtask



task SBOX();


PIM_Command(32'd84148864);
PIM_Command(32'd84345217);
PIM_Command(32'd84345986);
PIM_Command(32'd84345475);
PIM_Command(32'd84280725);
PIM_Command(32'd93651076);
PIM_Command(32'd92537989);
PIM_Command(32'd92373126);
PIM_Command(32'd92538759);
PIM_Command(32'd92537224);
PIM_Command(32'd92832649);
PIM_Command(32'd84117142);
PIM_Command(32'd93717130);
PIM_Command(32'd93718155);
PIM_Command(32'd92930188);
PIM_Command(32'd92968333);
PIM_Command(32'd93029006);
PIM_Command(32'd83922575);
PIM_Command(32'd93163152);
PIM_Command(32'd93160337);
PIM_Command(32'd93687442);
PIM_Command(32'd92377747);
PIM_Command(32'd84382356);
PIM_Command(32'd75926167);
PIM_Command(32'd76123288);
PIM_Command(32'd93886361);
PIM_Command(32'd75825306);
PIM_Command(32'd94017435);
PIM_Command(32'd75600540);
PIM_Command(32'd76055709);
PIM_Command(32'd94215326);
PIM_Command(32'd75992991);
PIM_Command(32'd94346400);
PIM_Command(32'd75665057);
PIM_Command(32'd75534498);
PIM_Command(32'd94544291);
PIM_Command(32'd75730340);
PIM_Command(32'd94675365);
PIM_Command(32'd93948838);
PIM_Command(32'd94086567);
PIM_Command(32'd94282664);
PIM_Command(32'd94414249);
PIM_Command(32'd94806954);
PIM_Command(32'd94867883);
PIM_Command(32'd94933932);
PIM_Command(32'd94999725);
PIM_Command(32'd95071150);
PIM_Command(32'd78294191);
PIM_Command(32'd95268784);
PIM_Command(32'd78557361);
PIM_Command(32'd95529906);
PIM_Command(32'd95202739);
PIM_Command(32'd95137716);
PIM_Command(32'd78951349);
PIM_Command(32'd95792566);
PIM_Command(32'd95205047);
PIM_Command(32'd95467192);
PIM_Command(32'd78493881);
PIM_Command(32'd96057274);
PIM_Command(32'd95467963);
PIM_Command(32'd78822332);
PIM_Command(32'd95337661);
PIM_Command(32'd96320190);
PIM_Command(32'd95598271);
PIM_Command(32'd95600064);
PIM_Command(32'd95861441);
PIM_Command(32'd96452290);
PIM_Command(32'd79792835);
PIM_Command(32'd79334596);
PIM_Command(32'd79036613);
PIM_Command(32'd79729350);
PIM_Command(32'd79529159);
PIM_Command(32'd78811080);
PIM_Command(32'd79662793);
PIM_Command(32'd79859914);
PIM_Command(32'd79597003);
PIM_Command(32'd79791820);
PIM_Command(32'd79333837);
PIM_Command(32'd79070670);
PIM_Command(32'd79725007);
PIM_Command(32'd79530192);
PIM_Command(32'd78809041);
PIM_Command(32'd79659730);
PIM_Command(32'd79855827);
PIM_Command(32'd79594452);
PIM_Command(32'd97702869);
PIM_Command(32'd97375702);
PIM_Command(32'd97310423);
PIM_Command(32'd96716248);
PIM_Command(32'd96781273);
PIM_Command(32'd96913370);
PIM_Command(32'd97507547);
PIM_Command(32'd97180380);
PIM_Command(32'd97246173);
PIM_Command(32'd98360798);
PIM_Command(32'd98228703);
PIM_Command(32'd96913632);
PIM_Command(32'd97572321);
PIM_Command(32'd98099426);
PIM_Command(32'd98033412);
PIM_Command(32'd97115363);
PIM_Command(32'd97640164);
PIM_Command(32'd98689765);
PIM_Command(32'd298837248);
PIM_Command(32'd97706982);
PIM_Command(32'd97963751);
PIM_Command(32'd98034439);
PIM_Command(32'd299820289);
PIM_Command(32'd98698243);
PIM_Command(32'd285532934);
PIM_Command(32'd98887400);
PIM_Command(32'd300471301);
PIM_Command(32'd99083266);
PIM_Command(32'd84675200);
PIM_Command(32'd84871553);
PIM_Command(32'd84872322);
PIM_Command(32'd84871811);
PIM_Command(32'd84807061);
PIM_Command(32'd93653124);
PIM_Command(32'd92540037);
PIM_Command(32'd92373126);
PIM_Command(32'd92540807);
PIM_Command(32'd92539272);
PIM_Command(32'd92832649);
PIM_Command(32'd84641430);
PIM_Command(32'd93719178);
PIM_Command(32'd93720203);
PIM_Command(32'd92932236);
PIM_Command(32'd92968333);
PIM_Command(32'd93029006);
PIM_Command(32'd84446863);
PIM_Command(32'd93163152);
PIM_Command(32'd93160337);
PIM_Command(32'd93687442);
PIM_Command(32'd92377747);
PIM_Command(32'd84906644);
PIM_Command(32'd75926167);
PIM_Command(32'd76123288);
PIM_Command(32'd93886361);
PIM_Command(32'd75827354);
PIM_Command(32'd94017435);
PIM_Command(32'd75600540);
PIM_Command(32'd76055709);
PIM_Command(32'd94215326);
PIM_Command(32'd75992991);
PIM_Command(32'd94346400);
PIM_Command(32'd75665057);
PIM_Command(32'd75534498);
PIM_Command(32'd94544291);
PIM_Command(32'd75730340);
PIM_Command(32'd94675365);
PIM_Command(32'd93948838);
PIM_Command(32'd94086567);
PIM_Command(32'd94282664);
PIM_Command(32'd94414249);
PIM_Command(32'd94806954);
PIM_Command(32'd94867883);
PIM_Command(32'd94933932);
PIM_Command(32'd94999725);
PIM_Command(32'd95071150);
PIM_Command(32'd78294191);
PIM_Command(32'd95268784);
PIM_Command(32'd78557361);
PIM_Command(32'd95529906);
PIM_Command(32'd95202739);
PIM_Command(32'd95137716);
PIM_Command(32'd78951349);
PIM_Command(32'd95792566);
PIM_Command(32'd95205047);
PIM_Command(32'd95467192);
PIM_Command(32'd78493881);
PIM_Command(32'd96057274);
PIM_Command(32'd95467963);
PIM_Command(32'd78822332);
PIM_Command(32'd95337661);
PIM_Command(32'd96320190);
PIM_Command(32'd95598271);
PIM_Command(32'd95600064);
PIM_Command(32'd95861441);
PIM_Command(32'd96452290);
PIM_Command(32'd79792835);
PIM_Command(32'd79334596);
PIM_Command(32'd79038661);
PIM_Command(32'd79729350);
PIM_Command(32'd79529159);
PIM_Command(32'd78811080);
PIM_Command(32'd79662793);
PIM_Command(32'd79859914);
PIM_Command(32'd79597003);
PIM_Command(32'd79791820);
PIM_Command(32'd79333837);
PIM_Command(32'd79070670);
PIM_Command(32'd79725007);
PIM_Command(32'd79530192);
PIM_Command(32'd78809041);
PIM_Command(32'd79659730);
PIM_Command(32'd79855827);
PIM_Command(32'd79594452);
PIM_Command(32'd97702869);
PIM_Command(32'd97375702);
PIM_Command(32'd97310423);
PIM_Command(32'd96716248);
PIM_Command(32'd96781273);
PIM_Command(32'd96913370);
PIM_Command(32'd97507547);
PIM_Command(32'd97180380);
PIM_Command(32'd97246173);
PIM_Command(32'd98360798);
PIM_Command(32'd98228703);
PIM_Command(32'd96913632);
PIM_Command(32'd97572321);
PIM_Command(32'd98099426);
PIM_Command(32'd98033420);
PIM_Command(32'd97115363);
PIM_Command(32'd97640164);
PIM_Command(32'd98689765);
PIM_Command(32'd298837256);
PIM_Command(32'd97706982);
PIM_Command(32'd97963751);
PIM_Command(32'd98034447);
PIM_Command(32'd299820297);
PIM_Command(32'd98700299);
PIM_Command(32'd286057230);
PIM_Command(32'd98887400);
PIM_Command(32'd300471309);
PIM_Command(32'd99083274);
PIM_Command(32'd85201536);
PIM_Command(32'd85397889);
PIM_Command(32'd85398658);
PIM_Command(32'd85398147);
PIM_Command(32'd85333397);
PIM_Command(32'd93655172);
PIM_Command(32'd92542085);
PIM_Command(32'd92373126);
PIM_Command(32'd92542855);
PIM_Command(32'd92541320);
PIM_Command(32'd92832649);
PIM_Command(32'd85165718);
PIM_Command(32'd93721226);
PIM_Command(32'd93722251);
PIM_Command(32'd92934284);
PIM_Command(32'd92968333);
PIM_Command(32'd93029006);
PIM_Command(32'd84971151);
PIM_Command(32'd93163152);
PIM_Command(32'd93160337);
PIM_Command(32'd93687442);
PIM_Command(32'd92377747);
PIM_Command(32'd85430932);
PIM_Command(32'd75926167);
PIM_Command(32'd76123288);
PIM_Command(32'd93886361);
PIM_Command(32'd75829402);
PIM_Command(32'd94017435);
PIM_Command(32'd75600540);
PIM_Command(32'd76055709);
PIM_Command(32'd94215326);
PIM_Command(32'd75992991);
PIM_Command(32'd94346400);
PIM_Command(32'd75665057);
PIM_Command(32'd75534498);
PIM_Command(32'd94544291);
PIM_Command(32'd75730340);
PIM_Command(32'd94675365);
PIM_Command(32'd93948838);
PIM_Command(32'd94086567);
PIM_Command(32'd94282664);
PIM_Command(32'd94414249);
PIM_Command(32'd94806954);
PIM_Command(32'd94867883);
PIM_Command(32'd94933932);
PIM_Command(32'd94999725);
PIM_Command(32'd95071150);
PIM_Command(32'd78294191);
PIM_Command(32'd95268784);
PIM_Command(32'd78557361);
PIM_Command(32'd95529906);
PIM_Command(32'd95202739);
PIM_Command(32'd95137716);
PIM_Command(32'd78951349);
PIM_Command(32'd95792566);
PIM_Command(32'd95205047);
PIM_Command(32'd95467192);
PIM_Command(32'd78493881);
PIM_Command(32'd96057274);
PIM_Command(32'd95467963);
PIM_Command(32'd78822332);
PIM_Command(32'd95337661);
PIM_Command(32'd96320190);
PIM_Command(32'd95598271);
PIM_Command(32'd95600064);
PIM_Command(32'd95861441);
PIM_Command(32'd96452290);
PIM_Command(32'd79792835);
PIM_Command(32'd79334596);
PIM_Command(32'd79040709);
PIM_Command(32'd79729350);
PIM_Command(32'd79529159);
PIM_Command(32'd78811080);
PIM_Command(32'd79662793);
PIM_Command(32'd79859914);
PIM_Command(32'd79597003);
PIM_Command(32'd79791820);
PIM_Command(32'd79333837);
PIM_Command(32'd79070670);
PIM_Command(32'd79725007);
PIM_Command(32'd79530192);
PIM_Command(32'd78809041);
PIM_Command(32'd79659730);
PIM_Command(32'd79855827);
PIM_Command(32'd79594452);
PIM_Command(32'd97702869);
PIM_Command(32'd97375702);
PIM_Command(32'd97310423);
PIM_Command(32'd96716248);
PIM_Command(32'd96781273);
PIM_Command(32'd96913370);
PIM_Command(32'd97507547);
PIM_Command(32'd97180380);
PIM_Command(32'd97246173);
PIM_Command(32'd98360798);
PIM_Command(32'd98228703);
PIM_Command(32'd96913632);
PIM_Command(32'd97572321);
PIM_Command(32'd98099426);
PIM_Command(32'd98033428);
PIM_Command(32'd97115363);
PIM_Command(32'd97640164);
PIM_Command(32'd98689765);
PIM_Command(32'd298837264);
PIM_Command(32'd97706982);
PIM_Command(32'd97963751);
PIM_Command(32'd98034455);
PIM_Command(32'd299820305);
PIM_Command(32'd98702355);
PIM_Command(32'd286581526);
PIM_Command(32'd98887400);
PIM_Command(32'd300471317);
PIM_Command(32'd99083282);
PIM_Command(32'd85727872);
PIM_Command(32'd85924225);
PIM_Command(32'd85924994);
PIM_Command(32'd85924483);
PIM_Command(32'd85859733);
PIM_Command(32'd93657220);
PIM_Command(32'd92544133);
PIM_Command(32'd92373126);
PIM_Command(32'd92544903);
PIM_Command(32'd92543368);
PIM_Command(32'd92832649);
PIM_Command(32'd85690006);
PIM_Command(32'd93723274);
PIM_Command(32'd93724299);
PIM_Command(32'd92936332);
PIM_Command(32'd92968333);
PIM_Command(32'd93029006);
PIM_Command(32'd85495439);
PIM_Command(32'd93163152);
PIM_Command(32'd93160337);
PIM_Command(32'd93687442);
PIM_Command(32'd92377747);
PIM_Command(32'd85955220);
PIM_Command(32'd75926167);
PIM_Command(32'd76123288);
PIM_Command(32'd93886361);
PIM_Command(32'd75831450);
PIM_Command(32'd94017435);
PIM_Command(32'd75600540);
PIM_Command(32'd76055709);
PIM_Command(32'd94215326);
PIM_Command(32'd75992991);
PIM_Command(32'd94346400);
PIM_Command(32'd75665057);
PIM_Command(32'd75534498);
PIM_Command(32'd94544291);
PIM_Command(32'd75730340);
PIM_Command(32'd94675365);
PIM_Command(32'd93948838);
PIM_Command(32'd94086567);
PIM_Command(32'd94282664);
PIM_Command(32'd94414249);
PIM_Command(32'd94806954);
PIM_Command(32'd94867883);
PIM_Command(32'd94933932);
PIM_Command(32'd94999725);
PIM_Command(32'd95071150);
PIM_Command(32'd78294191);
PIM_Command(32'd95268784);
PIM_Command(32'd78557361);
PIM_Command(32'd95529906);
PIM_Command(32'd95202739);
PIM_Command(32'd95137716);
PIM_Command(32'd78951349);
PIM_Command(32'd95792566);
PIM_Command(32'd95205047);
PIM_Command(32'd95467192);
PIM_Command(32'd78493881);
PIM_Command(32'd96057274);
PIM_Command(32'd95467963);
PIM_Command(32'd78822332);
PIM_Command(32'd95337661);
PIM_Command(32'd96320190);
PIM_Command(32'd95598271);
PIM_Command(32'd95600064);
PIM_Command(32'd95861441);
PIM_Command(32'd96452290);
PIM_Command(32'd79792835);
PIM_Command(32'd79334596);
PIM_Command(32'd79042757);
PIM_Command(32'd79729350);
PIM_Command(32'd79529159);
PIM_Command(32'd78811080);
PIM_Command(32'd79662793);
PIM_Command(32'd79859914);
PIM_Command(32'd79597003);
PIM_Command(32'd79791820);
PIM_Command(32'd79333837);
PIM_Command(32'd79070670);
PIM_Command(32'd79725007);
PIM_Command(32'd79530192);
PIM_Command(32'd78809041);
PIM_Command(32'd79659730);
PIM_Command(32'd79855827);
PIM_Command(32'd79594452);
PIM_Command(32'd97702869);
PIM_Command(32'd97375702);
PIM_Command(32'd97310423);
PIM_Command(32'd96716248);
PIM_Command(32'd96781273);
PIM_Command(32'd96913370);
PIM_Command(32'd97507547);
PIM_Command(32'd97180380);
PIM_Command(32'd97246173);
PIM_Command(32'd98360798);
PIM_Command(32'd98228703);
PIM_Command(32'd96913632);
PIM_Command(32'd97572321);
PIM_Command(32'd98099426);
PIM_Command(32'd98033436);
PIM_Command(32'd97115363);
PIM_Command(32'd97640164);
PIM_Command(32'd98689765);
PIM_Command(32'd298837272);
PIM_Command(32'd97706982);
PIM_Command(32'd97963751);
PIM_Command(32'd98034463);
PIM_Command(32'd299820313);
PIM_Command(32'd98704411);
PIM_Command(32'd287105822);
PIM_Command(32'd98887400);
PIM_Command(32'd300471325);
PIM_Command(32'd99083290);
PIM_Command(32'd86254208);
PIM_Command(32'd86450561);
PIM_Command(32'd86451330);
PIM_Command(32'd86450819);
PIM_Command(32'd86386069);
PIM_Command(32'd93659268);
PIM_Command(32'd92546181);
PIM_Command(32'd92373126);
PIM_Command(32'd92546951);
PIM_Command(32'd92545416);
PIM_Command(32'd92832649);
PIM_Command(32'd86214294);
PIM_Command(32'd93725322);
PIM_Command(32'd93726347);
PIM_Command(32'd92938380);
PIM_Command(32'd92968333);
PIM_Command(32'd93029006);
PIM_Command(32'd86019727);
PIM_Command(32'd93163152);
PIM_Command(32'd93160337);
PIM_Command(32'd93687442);
PIM_Command(32'd92377747);
PIM_Command(32'd86479508);
PIM_Command(32'd75926167);
PIM_Command(32'd76123288);
PIM_Command(32'd93886361);
PIM_Command(32'd75833498);
PIM_Command(32'd94017435);
PIM_Command(32'd75600540);
PIM_Command(32'd76055709);
PIM_Command(32'd94215326);
PIM_Command(32'd75992991);
PIM_Command(32'd94346400);
PIM_Command(32'd75665057);
PIM_Command(32'd75534498);
PIM_Command(32'd94544291);
PIM_Command(32'd75730340);
PIM_Command(32'd94675365);
PIM_Command(32'd93948838);
PIM_Command(32'd94086567);
PIM_Command(32'd94282664);
PIM_Command(32'd94414249);
PIM_Command(32'd94806954);
PIM_Command(32'd94867883);
PIM_Command(32'd94933932);
PIM_Command(32'd94999725);
PIM_Command(32'd95071150);
PIM_Command(32'd78294191);
PIM_Command(32'd95268784);
PIM_Command(32'd78557361);
PIM_Command(32'd95529906);
PIM_Command(32'd95202739);
PIM_Command(32'd95137716);
PIM_Command(32'd78951349);
PIM_Command(32'd95792566);
PIM_Command(32'd95205047);
PIM_Command(32'd95467192);
PIM_Command(32'd78493881);
PIM_Command(32'd96057274);
PIM_Command(32'd95467963);
PIM_Command(32'd78822332);
PIM_Command(32'd95337661);
PIM_Command(32'd96320190);
PIM_Command(32'd95598271);
PIM_Command(32'd95600064);
PIM_Command(32'd95861441);
PIM_Command(32'd96452290);
PIM_Command(32'd79792835);
PIM_Command(32'd79334596);
PIM_Command(32'd79044805);
PIM_Command(32'd79729350);
PIM_Command(32'd79529159);
PIM_Command(32'd78811080);
PIM_Command(32'd79662793);
PIM_Command(32'd79859914);
PIM_Command(32'd79597003);
PIM_Command(32'd79791820);
PIM_Command(32'd79333837);
PIM_Command(32'd79070670);
PIM_Command(32'd79725007);
PIM_Command(32'd79530192);
PIM_Command(32'd78809041);
PIM_Command(32'd79659730);
PIM_Command(32'd79855827);
PIM_Command(32'd79594452);
PIM_Command(32'd97702869);
PIM_Command(32'd97375702);
PIM_Command(32'd97310423);
PIM_Command(32'd96716248);
PIM_Command(32'd96781273);
PIM_Command(32'd96913370);
PIM_Command(32'd97507547);
PIM_Command(32'd97180380);
PIM_Command(32'd97246173);
PIM_Command(32'd98360798);
PIM_Command(32'd98228703);
PIM_Command(32'd96913632);
PIM_Command(32'd97572321);
PIM_Command(32'd98099426);
PIM_Command(32'd98033444);
PIM_Command(32'd97115363);
PIM_Command(32'd97640164);
PIM_Command(32'd98689765);
PIM_Command(32'd298837280);
PIM_Command(32'd97706982);
PIM_Command(32'd97963751);
PIM_Command(32'd98034471);
PIM_Command(32'd299820321);
PIM_Command(32'd98706467);
PIM_Command(32'd287630118);
PIM_Command(32'd98887400);
PIM_Command(32'd300471333);
PIM_Command(32'd99083298);
PIM_Command(32'd86780544);
PIM_Command(32'd86976897);
PIM_Command(32'd86977666);
PIM_Command(32'd86977155);
PIM_Command(32'd86912405);
PIM_Command(32'd93661316);
PIM_Command(32'd92548229);
PIM_Command(32'd92373126);
PIM_Command(32'd92548999);
PIM_Command(32'd92547464);
PIM_Command(32'd92832649);
PIM_Command(32'd86738582);
PIM_Command(32'd93727370);
PIM_Command(32'd93728395);
PIM_Command(32'd92940428);
PIM_Command(32'd92968333);
PIM_Command(32'd93029006);
PIM_Command(32'd86544015);
PIM_Command(32'd93163152);
PIM_Command(32'd93160337);
PIM_Command(32'd93687442);
PIM_Command(32'd92377747);
PIM_Command(32'd87003796);
PIM_Command(32'd75926167);
PIM_Command(32'd76123288);
PIM_Command(32'd93886361);
PIM_Command(32'd75835546);
PIM_Command(32'd94017435);
PIM_Command(32'd75600540);
PIM_Command(32'd76055709);
PIM_Command(32'd94215326);
PIM_Command(32'd75992991);
PIM_Command(32'd94346400);
PIM_Command(32'd75665057);
PIM_Command(32'd75534498);
PIM_Command(32'd94544291);
PIM_Command(32'd75730340);
PIM_Command(32'd94675365);
PIM_Command(32'd93948838);
PIM_Command(32'd94086567);
PIM_Command(32'd94282664);
PIM_Command(32'd94414249);
PIM_Command(32'd94806954);
PIM_Command(32'd94867883);
PIM_Command(32'd94933932);
PIM_Command(32'd94999725);
PIM_Command(32'd95071150);
PIM_Command(32'd78294191);
PIM_Command(32'd95268784);
PIM_Command(32'd78557361);
PIM_Command(32'd95529906);
PIM_Command(32'd95202739);
PIM_Command(32'd95137716);
PIM_Command(32'd78951349);
PIM_Command(32'd95792566);
PIM_Command(32'd95205047);
PIM_Command(32'd95467192);
PIM_Command(32'd78493881);
PIM_Command(32'd96057274);
PIM_Command(32'd95467963);
PIM_Command(32'd78822332);
PIM_Command(32'd95337661);
PIM_Command(32'd96320190);
PIM_Command(32'd95598271);
PIM_Command(32'd95600064);
PIM_Command(32'd95861441);
PIM_Command(32'd96452290);
PIM_Command(32'd79792835);
PIM_Command(32'd79334596);
PIM_Command(32'd79046853);
PIM_Command(32'd79729350);
PIM_Command(32'd79529159);
PIM_Command(32'd78811080);
PIM_Command(32'd79662793);
PIM_Command(32'd79859914);
PIM_Command(32'd79597003);
PIM_Command(32'd79791820);
PIM_Command(32'd79333837);
PIM_Command(32'd79070670);
PIM_Command(32'd79725007);
PIM_Command(32'd79530192);
PIM_Command(32'd78809041);
PIM_Command(32'd79659730);
PIM_Command(32'd79855827);
PIM_Command(32'd79594452);
PIM_Command(32'd97702869);
PIM_Command(32'd97375702);
PIM_Command(32'd97310423);
PIM_Command(32'd96716248);
PIM_Command(32'd96781273);
PIM_Command(32'd96913370);
PIM_Command(32'd97507547);
PIM_Command(32'd97180380);
PIM_Command(32'd97246173);
PIM_Command(32'd98360798);
PIM_Command(32'd98228703);
PIM_Command(32'd96913632);
PIM_Command(32'd97572321);
PIM_Command(32'd98099426);
PIM_Command(32'd98033452);
PIM_Command(32'd97115363);
PIM_Command(32'd97640164);
PIM_Command(32'd98689765);
PIM_Command(32'd298837288);
PIM_Command(32'd97706982);
PIM_Command(32'd97963751);
PIM_Command(32'd98034479);
PIM_Command(32'd299820329);
PIM_Command(32'd98708523);
PIM_Command(32'd288154414);
PIM_Command(32'd98887400);
PIM_Command(32'd300471341);
PIM_Command(32'd99083306);
PIM_Command(32'd87306880);
PIM_Command(32'd87503233);
PIM_Command(32'd87504002);
PIM_Command(32'd87503491);
PIM_Command(32'd87438741);
PIM_Command(32'd93663364);
PIM_Command(32'd92550277);
PIM_Command(32'd92373126);
PIM_Command(32'd92551047);
PIM_Command(32'd92549512);
PIM_Command(32'd92832649);
PIM_Command(32'd87262870);
PIM_Command(32'd93729418);
PIM_Command(32'd93730443);
PIM_Command(32'd92942476);
PIM_Command(32'd92968333);
PIM_Command(32'd93029006);
PIM_Command(32'd87068303);
PIM_Command(32'd93163152);
PIM_Command(32'd93160337);
PIM_Command(32'd93687442);
PIM_Command(32'd92377747);
PIM_Command(32'd87528084);
PIM_Command(32'd75926167);
PIM_Command(32'd76123288);
PIM_Command(32'd93886361);
PIM_Command(32'd75837594);
PIM_Command(32'd94017435);
PIM_Command(32'd75600540);
PIM_Command(32'd76055709);
PIM_Command(32'd94215326);
PIM_Command(32'd75992991);
PIM_Command(32'd94346400);
PIM_Command(32'd75665057);
PIM_Command(32'd75534498);
PIM_Command(32'd94544291);
PIM_Command(32'd75730340);
PIM_Command(32'd94675365);
PIM_Command(32'd93948838);
PIM_Command(32'd94086567);
PIM_Command(32'd94282664);
PIM_Command(32'd94414249);
PIM_Command(32'd94806954);
PIM_Command(32'd94867883);
PIM_Command(32'd94933932);
PIM_Command(32'd94999725);
PIM_Command(32'd95071150);
PIM_Command(32'd78294191);
PIM_Command(32'd95268784);
PIM_Command(32'd78557361);
PIM_Command(32'd95529906);
PIM_Command(32'd95202739);
PIM_Command(32'd95137716);
PIM_Command(32'd78951349);
PIM_Command(32'd95792566);
PIM_Command(32'd95205047);
PIM_Command(32'd95467192);
PIM_Command(32'd78493881);
PIM_Command(32'd96057274);
PIM_Command(32'd95467963);
PIM_Command(32'd78822332);
PIM_Command(32'd95337661);
PIM_Command(32'd96320190);
PIM_Command(32'd95598271);
PIM_Command(32'd95600064);
PIM_Command(32'd95861441);
PIM_Command(32'd96452290);
PIM_Command(32'd79792835);
PIM_Command(32'd79334596);
PIM_Command(32'd79048901);
PIM_Command(32'd79729350);
PIM_Command(32'd79529159);
PIM_Command(32'd78811080);
PIM_Command(32'd79662793);
PIM_Command(32'd79859914);
PIM_Command(32'd79597003);
PIM_Command(32'd79791820);
PIM_Command(32'd79333837);
PIM_Command(32'd79070670);
PIM_Command(32'd79725007);
PIM_Command(32'd79530192);
PIM_Command(32'd78809041);
PIM_Command(32'd79659730);
PIM_Command(32'd79855827);
PIM_Command(32'd79594452);
PIM_Command(32'd97702869);
PIM_Command(32'd97375702);
PIM_Command(32'd97310423);
PIM_Command(32'd96716248);
PIM_Command(32'd96781273);
PIM_Command(32'd96913370);
PIM_Command(32'd97507547);
PIM_Command(32'd97180380);
PIM_Command(32'd97246173);
PIM_Command(32'd98360798);
PIM_Command(32'd98228703);
PIM_Command(32'd96913632);
PIM_Command(32'd97572321);
PIM_Command(32'd98099426);
PIM_Command(32'd98033460);
PIM_Command(32'd97115363);
PIM_Command(32'd97640164);
PIM_Command(32'd98689765);
PIM_Command(32'd298837296);
PIM_Command(32'd97706982);
PIM_Command(32'd97963751);
PIM_Command(32'd98034487);
PIM_Command(32'd299820337);
PIM_Command(32'd98710579);
PIM_Command(32'd288678710);
PIM_Command(32'd98887400);
PIM_Command(32'd300471349);
PIM_Command(32'd99083314);
PIM_Command(32'd87833216);
PIM_Command(32'd88029569);
PIM_Command(32'd88030338);
PIM_Command(32'd88029827);
PIM_Command(32'd87965077);
PIM_Command(32'd93665412);
PIM_Command(32'd92552325);
PIM_Command(32'd92373126);
PIM_Command(32'd92553095);
PIM_Command(32'd92551560);
PIM_Command(32'd92832649);
PIM_Command(32'd87787158);
PIM_Command(32'd93731466);
PIM_Command(32'd93732491);
PIM_Command(32'd92944524);
PIM_Command(32'd92968333);
PIM_Command(32'd93029006);
PIM_Command(32'd87592591);
PIM_Command(32'd93163152);
PIM_Command(32'd93160337);
PIM_Command(32'd93687442);
PIM_Command(32'd92377747);
PIM_Command(32'd88052372);
PIM_Command(32'd75926167);
PIM_Command(32'd76123288);
PIM_Command(32'd93886361);
PIM_Command(32'd75839642);
PIM_Command(32'd94017435);
PIM_Command(32'd75600540);
PIM_Command(32'd76055709);
PIM_Command(32'd94215326);
PIM_Command(32'd75992991);
PIM_Command(32'd94346400);
PIM_Command(32'd75665057);
PIM_Command(32'd75534498);
PIM_Command(32'd94544291);
PIM_Command(32'd75730340);
PIM_Command(32'd94675365);
PIM_Command(32'd93948838);
PIM_Command(32'd94086567);
PIM_Command(32'd94282664);
PIM_Command(32'd94414249);
PIM_Command(32'd94806954);
PIM_Command(32'd94867883);
PIM_Command(32'd94933932);
PIM_Command(32'd94999725);
PIM_Command(32'd95071150);
PIM_Command(32'd78294191);
PIM_Command(32'd95268784);
PIM_Command(32'd78557361);
PIM_Command(32'd95529906);
PIM_Command(32'd95202739);
PIM_Command(32'd95137716);
PIM_Command(32'd78951349);
PIM_Command(32'd95792566);
PIM_Command(32'd95205047);
PIM_Command(32'd95467192);
PIM_Command(32'd78493881);
PIM_Command(32'd96057274);
PIM_Command(32'd95467963);
PIM_Command(32'd78822332);
PIM_Command(32'd95337661);
PIM_Command(32'd96320190);
PIM_Command(32'd95598271);
PIM_Command(32'd95600064);
PIM_Command(32'd95861441);
PIM_Command(32'd96452290);
PIM_Command(32'd79792835);
PIM_Command(32'd79334596);
PIM_Command(32'd79050949);
PIM_Command(32'd79729350);
PIM_Command(32'd79529159);
PIM_Command(32'd78811080);
PIM_Command(32'd79662793);
PIM_Command(32'd79859914);
PIM_Command(32'd79597003);
PIM_Command(32'd79791820);
PIM_Command(32'd79333837);
PIM_Command(32'd79070670);
PIM_Command(32'd79725007);
PIM_Command(32'd79530192);
PIM_Command(32'd78809041);
PIM_Command(32'd79659730);
PIM_Command(32'd79855827);
PIM_Command(32'd79594452);
PIM_Command(32'd97702869);
PIM_Command(32'd97375702);
PIM_Command(32'd97310423);
PIM_Command(32'd96716248);
PIM_Command(32'd96781273);
PIM_Command(32'd96913370);
PIM_Command(32'd97507547);
PIM_Command(32'd97180380);
PIM_Command(32'd97246173);
PIM_Command(32'd98360798);
PIM_Command(32'd98228703);
PIM_Command(32'd96913632);
PIM_Command(32'd97572321);
PIM_Command(32'd98099426);
PIM_Command(32'd98033468);
PIM_Command(32'd97115363);
PIM_Command(32'd97640164);
PIM_Command(32'd98689765);
PIM_Command(32'd298837304);
PIM_Command(32'd97706982);
PIM_Command(32'd97963751);
PIM_Command(32'd98034495);
PIM_Command(32'd299820345);
PIM_Command(32'd98712635);
PIM_Command(32'd289203006);
PIM_Command(32'd98887400);
PIM_Command(32'd300471357);
PIM_Command(32'd99083322);
PIM_Command(32'd88359552);
PIM_Command(32'd88555905);
PIM_Command(32'd88556674);
PIM_Command(32'd88556163);
PIM_Command(32'd88491413);
PIM_Command(32'd93667460);
PIM_Command(32'd92554373);
PIM_Command(32'd92373126);
PIM_Command(32'd92555143);
PIM_Command(32'd92553608);
PIM_Command(32'd92832649);
PIM_Command(32'd88311446);
PIM_Command(32'd93733514);
PIM_Command(32'd93734539);
PIM_Command(32'd92946572);
PIM_Command(32'd92968333);
PIM_Command(32'd93029006);
PIM_Command(32'd88116879);
PIM_Command(32'd93163152);
PIM_Command(32'd93160337);
PIM_Command(32'd93687442);
PIM_Command(32'd92377747);
PIM_Command(32'd88576660);
PIM_Command(32'd75926167);
PIM_Command(32'd76123288);
PIM_Command(32'd93886361);
PIM_Command(32'd75841690);
PIM_Command(32'd94017435);
PIM_Command(32'd75600540);
PIM_Command(32'd76055709);
PIM_Command(32'd94215326);
PIM_Command(32'd75992991);
PIM_Command(32'd94346400);
PIM_Command(32'd75665057);
PIM_Command(32'd75534498);
PIM_Command(32'd94544291);
PIM_Command(32'd75730340);
PIM_Command(32'd94675365);
PIM_Command(32'd93948838);
PIM_Command(32'd94086567);
PIM_Command(32'd94282664);
PIM_Command(32'd94414249);
PIM_Command(32'd94806954);
PIM_Command(32'd94867883);
PIM_Command(32'd94933932);
PIM_Command(32'd94999725);
PIM_Command(32'd95071150);
PIM_Command(32'd78294191);
PIM_Command(32'd95268784);
PIM_Command(32'd78557361);
PIM_Command(32'd95529906);
PIM_Command(32'd95202739);
PIM_Command(32'd95137716);
PIM_Command(32'd78951349);
PIM_Command(32'd95792566);
PIM_Command(32'd95205047);
PIM_Command(32'd95467192);
PIM_Command(32'd78493881);
PIM_Command(32'd96057274);
PIM_Command(32'd95467963);
PIM_Command(32'd78822332);
PIM_Command(32'd95337661);
PIM_Command(32'd96320190);
PIM_Command(32'd95598271);
PIM_Command(32'd95600064);
PIM_Command(32'd95861441);
PIM_Command(32'd96452290);
PIM_Command(32'd79792835);
PIM_Command(32'd79334596);
PIM_Command(32'd79052997);
PIM_Command(32'd79729350);
PIM_Command(32'd79529159);
PIM_Command(32'd78811080);
PIM_Command(32'd79662793);
PIM_Command(32'd79859914);
PIM_Command(32'd79597003);
PIM_Command(32'd79791820);
PIM_Command(32'd79333837);
PIM_Command(32'd79070670);
PIM_Command(32'd79725007);
PIM_Command(32'd79530192);
PIM_Command(32'd78809041);
PIM_Command(32'd79659730);
PIM_Command(32'd79855827);
PIM_Command(32'd79594452);
PIM_Command(32'd97702869);
PIM_Command(32'd97375702);
PIM_Command(32'd97310423);
PIM_Command(32'd96716248);
PIM_Command(32'd96781273);
PIM_Command(32'd96913370);
PIM_Command(32'd97507547);
PIM_Command(32'd97180380);
PIM_Command(32'd97246173);
PIM_Command(32'd98360798);
PIM_Command(32'd98228703);
PIM_Command(32'd96913632);
PIM_Command(32'd97572321);
PIM_Command(32'd98099426);
PIM_Command(32'd98033476);
PIM_Command(32'd97115363);
PIM_Command(32'd97640164);
PIM_Command(32'd98689765);
PIM_Command(32'd298837312);
PIM_Command(32'd97706982);
PIM_Command(32'd97963751);
PIM_Command(32'd98034503);
PIM_Command(32'd299820353);
PIM_Command(32'd98714691);
PIM_Command(32'd289727302);
PIM_Command(32'd98887400);
PIM_Command(32'd300471365);
PIM_Command(32'd99083330);
PIM_Command(32'd88885888);
PIM_Command(32'd89082241);
PIM_Command(32'd89083010);
PIM_Command(32'd89082499);
PIM_Command(32'd89017749);
PIM_Command(32'd93669508);
PIM_Command(32'd92556421);
PIM_Command(32'd92373126);
PIM_Command(32'd92557191);
PIM_Command(32'd92555656);
PIM_Command(32'd92832649);
PIM_Command(32'd88835734);
PIM_Command(32'd93735562);
PIM_Command(32'd93736587);
PIM_Command(32'd92948620);
PIM_Command(32'd92968333);
PIM_Command(32'd93029006);
PIM_Command(32'd88641167);
PIM_Command(32'd93163152);
PIM_Command(32'd93160337);
PIM_Command(32'd93687442);
PIM_Command(32'd92377747);
PIM_Command(32'd89100948);
PIM_Command(32'd75926167);
PIM_Command(32'd76123288);
PIM_Command(32'd93886361);
PIM_Command(32'd75843738);
PIM_Command(32'd94017435);
PIM_Command(32'd75600540);
PIM_Command(32'd76055709);
PIM_Command(32'd94215326);
PIM_Command(32'd75992991);
PIM_Command(32'd94346400);
PIM_Command(32'd75665057);
PIM_Command(32'd75534498);
PIM_Command(32'd94544291);
PIM_Command(32'd75730340);
PIM_Command(32'd94675365);
PIM_Command(32'd93948838);
PIM_Command(32'd94086567);
PIM_Command(32'd94282664);
PIM_Command(32'd94414249);
PIM_Command(32'd94806954);
PIM_Command(32'd94867883);
PIM_Command(32'd94933932);
PIM_Command(32'd94999725);
PIM_Command(32'd95071150);
PIM_Command(32'd78294191);
PIM_Command(32'd95268784);
PIM_Command(32'd78557361);
PIM_Command(32'd95529906);
PIM_Command(32'd95202739);
PIM_Command(32'd95137716);
PIM_Command(32'd78951349);
PIM_Command(32'd95792566);
PIM_Command(32'd95205047);
PIM_Command(32'd95467192);
PIM_Command(32'd78493881);
PIM_Command(32'd96057274);
PIM_Command(32'd95467963);
PIM_Command(32'd78822332);
PIM_Command(32'd95337661);
PIM_Command(32'd96320190);
PIM_Command(32'd95598271);
PIM_Command(32'd95600064);
PIM_Command(32'd95861441);
PIM_Command(32'd96452290);
PIM_Command(32'd79792835);
PIM_Command(32'd79334596);
PIM_Command(32'd79055045);
PIM_Command(32'd79729350);
PIM_Command(32'd79529159);
PIM_Command(32'd78811080);
PIM_Command(32'd79662793);
PIM_Command(32'd79859914);
PIM_Command(32'd79597003);
PIM_Command(32'd79791820);
PIM_Command(32'd79333837);
PIM_Command(32'd79070670);
PIM_Command(32'd79725007);
PIM_Command(32'd79530192);
PIM_Command(32'd78809041);
PIM_Command(32'd79659730);
PIM_Command(32'd79855827);
PIM_Command(32'd79594452);
PIM_Command(32'd97702869);
PIM_Command(32'd97375702);
PIM_Command(32'd97310423);
PIM_Command(32'd96716248);
PIM_Command(32'd96781273);
PIM_Command(32'd96913370);
PIM_Command(32'd97507547);
PIM_Command(32'd97180380);
PIM_Command(32'd97246173);
PIM_Command(32'd98360798);
PIM_Command(32'd98228703);
PIM_Command(32'd96913632);
PIM_Command(32'd97572321);
PIM_Command(32'd98099426);
PIM_Command(32'd98033484);
PIM_Command(32'd97115363);
PIM_Command(32'd97640164);
PIM_Command(32'd98689765);
PIM_Command(32'd298837320);
PIM_Command(32'd97706982);
PIM_Command(32'd97963751);
PIM_Command(32'd98034511);
PIM_Command(32'd299820361);
PIM_Command(32'd98716747);
PIM_Command(32'd290251598);
PIM_Command(32'd98887400);
PIM_Command(32'd300471373);
PIM_Command(32'd99083338);
PIM_Command(32'd89412224);
PIM_Command(32'd89608577);
PIM_Command(32'd89609346);
PIM_Command(32'd89608835);
PIM_Command(32'd89544085);
PIM_Command(32'd93671556);
PIM_Command(32'd92558469);
PIM_Command(32'd92373126);
PIM_Command(32'd92559239);
PIM_Command(32'd92557704);
PIM_Command(32'd92832649);
PIM_Command(32'd89360022);
PIM_Command(32'd93737610);
PIM_Command(32'd93738635);
PIM_Command(32'd92950668);
PIM_Command(32'd92968333);
PIM_Command(32'd93029006);
PIM_Command(32'd89165455);
PIM_Command(32'd93163152);
PIM_Command(32'd93160337);
PIM_Command(32'd93687442);
PIM_Command(32'd92377747);
PIM_Command(32'd89625236);
PIM_Command(32'd75926167);
PIM_Command(32'd76123288);
PIM_Command(32'd93886361);
PIM_Command(32'd75845786);
PIM_Command(32'd94017435);
PIM_Command(32'd75600540);
PIM_Command(32'd76055709);
PIM_Command(32'd94215326);
PIM_Command(32'd75992991);
PIM_Command(32'd94346400);
PIM_Command(32'd75665057);
PIM_Command(32'd75534498);
PIM_Command(32'd94544291);
PIM_Command(32'd75730340);
PIM_Command(32'd94675365);
PIM_Command(32'd93948838);
PIM_Command(32'd94086567);
PIM_Command(32'd94282664);
PIM_Command(32'd94414249);
PIM_Command(32'd94806954);
PIM_Command(32'd94867883);
PIM_Command(32'd94933932);
PIM_Command(32'd94999725);
PIM_Command(32'd95071150);
PIM_Command(32'd78294191);
PIM_Command(32'd95268784);
PIM_Command(32'd78557361);
PIM_Command(32'd95529906);
PIM_Command(32'd95202739);
PIM_Command(32'd95137716);
PIM_Command(32'd78951349);
PIM_Command(32'd95792566);
PIM_Command(32'd95205047);
PIM_Command(32'd95467192);
PIM_Command(32'd78493881);
PIM_Command(32'd96057274);
PIM_Command(32'd95467963);
PIM_Command(32'd78822332);
PIM_Command(32'd95337661);
PIM_Command(32'd96320190);
PIM_Command(32'd95598271);
PIM_Command(32'd95600064);
PIM_Command(32'd95861441);
PIM_Command(32'd96452290);
PIM_Command(32'd79792835);
PIM_Command(32'd79334596);
PIM_Command(32'd79057093);
PIM_Command(32'd79729350);
PIM_Command(32'd79529159);
PIM_Command(32'd78811080);
PIM_Command(32'd79662793);
PIM_Command(32'd79859914);
PIM_Command(32'd79597003);
PIM_Command(32'd79791820);
PIM_Command(32'd79333837);
PIM_Command(32'd79070670);
PIM_Command(32'd79725007);
PIM_Command(32'd79530192);
PIM_Command(32'd78809041);
PIM_Command(32'd79659730);
PIM_Command(32'd79855827);
PIM_Command(32'd79594452);
PIM_Command(32'd97702869);
PIM_Command(32'd97375702);
PIM_Command(32'd97310423);
PIM_Command(32'd96716248);
PIM_Command(32'd96781273);
PIM_Command(32'd96913370);
PIM_Command(32'd97507547);
PIM_Command(32'd97180380);
PIM_Command(32'd97246173);
PIM_Command(32'd98360798);
PIM_Command(32'd98228703);
PIM_Command(32'd96913632);
PIM_Command(32'd97572321);
PIM_Command(32'd98099426);
PIM_Command(32'd98033492);
PIM_Command(32'd97115363);
PIM_Command(32'd97640164);
PIM_Command(32'd98689765);
PIM_Command(32'd298837328);
PIM_Command(32'd97706982);
PIM_Command(32'd97963751);
PIM_Command(32'd98034519);
PIM_Command(32'd299820369);
PIM_Command(32'd98718803);
PIM_Command(32'd290775894);
PIM_Command(32'd98887400);
PIM_Command(32'd300471381);
PIM_Command(32'd99083346);
PIM_Command(32'd89938560);
PIM_Command(32'd90134913);
PIM_Command(32'd90135682);
PIM_Command(32'd90135171);
PIM_Command(32'd90070421);
PIM_Command(32'd93673604);
PIM_Command(32'd92560517);
PIM_Command(32'd92373126);
PIM_Command(32'd92561287);
PIM_Command(32'd92559752);
PIM_Command(32'd92832649);
PIM_Command(32'd89884310);
PIM_Command(32'd93739658);
PIM_Command(32'd93740683);
PIM_Command(32'd92952716);
PIM_Command(32'd92968333);
PIM_Command(32'd93029006);
PIM_Command(32'd89689743);
PIM_Command(32'd93163152);
PIM_Command(32'd93160337);
PIM_Command(32'd93687442);
PIM_Command(32'd92377747);
PIM_Command(32'd90149524);
PIM_Command(32'd75926167);
PIM_Command(32'd76123288);
PIM_Command(32'd93886361);
PIM_Command(32'd75847834);
PIM_Command(32'd94017435);
PIM_Command(32'd75600540);
PIM_Command(32'd76055709);
PIM_Command(32'd94215326);
PIM_Command(32'd75992991);
PIM_Command(32'd94346400);
PIM_Command(32'd75665057);
PIM_Command(32'd75534498);
PIM_Command(32'd94544291);
PIM_Command(32'd75730340);
PIM_Command(32'd94675365);
PIM_Command(32'd93948838);
PIM_Command(32'd94086567);
PIM_Command(32'd94282664);
PIM_Command(32'd94414249);
PIM_Command(32'd94806954);
PIM_Command(32'd94867883);
PIM_Command(32'd94933932);
PIM_Command(32'd94999725);
PIM_Command(32'd95071150);
PIM_Command(32'd78294191);
PIM_Command(32'd95268784);
PIM_Command(32'd78557361);
PIM_Command(32'd95529906);
PIM_Command(32'd95202739);
PIM_Command(32'd95137716);
PIM_Command(32'd78951349);
PIM_Command(32'd95792566);
PIM_Command(32'd95205047);
PIM_Command(32'd95467192);
PIM_Command(32'd78493881);
PIM_Command(32'd96057274);
PIM_Command(32'd95467963);
PIM_Command(32'd78822332);
PIM_Command(32'd95337661);
PIM_Command(32'd96320190);
PIM_Command(32'd95598271);
PIM_Command(32'd95600064);
PIM_Command(32'd95861441);
PIM_Command(32'd96452290);
PIM_Command(32'd79792835);
PIM_Command(32'd79334596);
PIM_Command(32'd79059141);
PIM_Command(32'd79729350);
PIM_Command(32'd79529159);
PIM_Command(32'd78811080);
PIM_Command(32'd79662793);
PIM_Command(32'd79859914);
PIM_Command(32'd79597003);
PIM_Command(32'd79791820);
PIM_Command(32'd79333837);
PIM_Command(32'd79070670);
PIM_Command(32'd79725007);
PIM_Command(32'd79530192);
PIM_Command(32'd78809041);
PIM_Command(32'd79659730);
PIM_Command(32'd79855827);
PIM_Command(32'd79594452);
PIM_Command(32'd97702869);
PIM_Command(32'd97375702);
PIM_Command(32'd97310423);
PIM_Command(32'd96716248);
PIM_Command(32'd96781273);
PIM_Command(32'd96913370);
PIM_Command(32'd97507547);
PIM_Command(32'd97180380);
PIM_Command(32'd97246173);
PIM_Command(32'd98360798);
PIM_Command(32'd98228703);
PIM_Command(32'd96913632);
PIM_Command(32'd97572321);
PIM_Command(32'd98099426);
PIM_Command(32'd98033500);
PIM_Command(32'd97115363);
PIM_Command(32'd97640164);
PIM_Command(32'd98689765);
PIM_Command(32'd298837336);
PIM_Command(32'd97706982);
PIM_Command(32'd97963751);
PIM_Command(32'd98034527);
PIM_Command(32'd299820377);
PIM_Command(32'd98720859);
PIM_Command(32'd291300190);
PIM_Command(32'd98887400);
PIM_Command(32'd300471389);
PIM_Command(32'd99083354);
PIM_Command(32'd90464896);
PIM_Command(32'd90661249);
PIM_Command(32'd90662018);
PIM_Command(32'd90661507);
PIM_Command(32'd90596757);
PIM_Command(32'd93675652);
PIM_Command(32'd92562565);
PIM_Command(32'd92373126);
PIM_Command(32'd92563335);
PIM_Command(32'd92561800);
PIM_Command(32'd92832649);
PIM_Command(32'd90408598);
PIM_Command(32'd93741706);
PIM_Command(32'd93742731);
PIM_Command(32'd92954764);
PIM_Command(32'd92968333);
PIM_Command(32'd93029006);
PIM_Command(32'd90214031);
PIM_Command(32'd93163152);
PIM_Command(32'd93160337);
PIM_Command(32'd93687442);
PIM_Command(32'd92377747);
PIM_Command(32'd90673812);
PIM_Command(32'd75926167);
PIM_Command(32'd76123288);
PIM_Command(32'd93886361);
PIM_Command(32'd75849882);
PIM_Command(32'd94017435);
PIM_Command(32'd75600540);
PIM_Command(32'd76055709);
PIM_Command(32'd94215326);
PIM_Command(32'd75992991);
PIM_Command(32'd94346400);
PIM_Command(32'd75665057);
PIM_Command(32'd75534498);
PIM_Command(32'd94544291);
PIM_Command(32'd75730340);
PIM_Command(32'd94675365);
PIM_Command(32'd93948838);
PIM_Command(32'd94086567);
PIM_Command(32'd94282664);
PIM_Command(32'd94414249);
PIM_Command(32'd94806954);
PIM_Command(32'd94867883);
PIM_Command(32'd94933932);
PIM_Command(32'd94999725);
PIM_Command(32'd95071150);
PIM_Command(32'd78294191);
PIM_Command(32'd95268784);
PIM_Command(32'd78557361);
PIM_Command(32'd95529906);
PIM_Command(32'd95202739);
PIM_Command(32'd95137716);
PIM_Command(32'd78951349);
PIM_Command(32'd95792566);
PIM_Command(32'd95205047);
PIM_Command(32'd95467192);
PIM_Command(32'd78493881);
PIM_Command(32'd96057274);
PIM_Command(32'd95467963);
PIM_Command(32'd78822332);
PIM_Command(32'd95337661);
PIM_Command(32'd96320190);
PIM_Command(32'd95598271);
PIM_Command(32'd95600064);
PIM_Command(32'd95861441);
PIM_Command(32'd96452290);
PIM_Command(32'd79792835);
PIM_Command(32'd79334596);
PIM_Command(32'd79061189);
PIM_Command(32'd79729350);
PIM_Command(32'd79529159);
PIM_Command(32'd78811080);
PIM_Command(32'd79662793);
PIM_Command(32'd79859914);
PIM_Command(32'd79597003);
PIM_Command(32'd79791820);
PIM_Command(32'd79333837);
PIM_Command(32'd79070670);
PIM_Command(32'd79725007);
PIM_Command(32'd79530192);
PIM_Command(32'd78809041);
PIM_Command(32'd79659730);
PIM_Command(32'd79855827);
PIM_Command(32'd79594452);
PIM_Command(32'd97702869);
PIM_Command(32'd97375702);
PIM_Command(32'd97310423);
PIM_Command(32'd96716248);
PIM_Command(32'd96781273);
PIM_Command(32'd96913370);
PIM_Command(32'd97507547);
PIM_Command(32'd97180380);
PIM_Command(32'd97246173);
PIM_Command(32'd98360798);
PIM_Command(32'd98228703);
PIM_Command(32'd96913632);
PIM_Command(32'd97572321);
PIM_Command(32'd98099426);
PIM_Command(32'd98033508);
PIM_Command(32'd97115363);
PIM_Command(32'd97640164);
PIM_Command(32'd98689765);
PIM_Command(32'd298837344);
PIM_Command(32'd97706982);
PIM_Command(32'd97963751);
PIM_Command(32'd98034535);
PIM_Command(32'd299820385);
PIM_Command(32'd98722915);
PIM_Command(32'd291824486);
PIM_Command(32'd98887400);
PIM_Command(32'd300471397);
PIM_Command(32'd99083362);
PIM_Command(32'd90991232);
PIM_Command(32'd91187585);
PIM_Command(32'd91188354);
PIM_Command(32'd91187843);
PIM_Command(32'd91123093);
PIM_Command(32'd93677700);
PIM_Command(32'd92564613);
PIM_Command(32'd92373126);
PIM_Command(32'd92565383);
PIM_Command(32'd92563848);
PIM_Command(32'd92832649);
PIM_Command(32'd90932886);
PIM_Command(32'd93743754);
PIM_Command(32'd93744779);
PIM_Command(32'd92956812);
PIM_Command(32'd92968333);
PIM_Command(32'd93029006);
PIM_Command(32'd90738319);
PIM_Command(32'd93163152);
PIM_Command(32'd93160337);
PIM_Command(32'd93687442);
PIM_Command(32'd92377747);
PIM_Command(32'd91198100);
PIM_Command(32'd75926167);
PIM_Command(32'd76123288);
PIM_Command(32'd93886361);
PIM_Command(32'd75851930);
PIM_Command(32'd94017435);
PIM_Command(32'd75600540);
PIM_Command(32'd76055709);
PIM_Command(32'd94215326);
PIM_Command(32'd75992991);
PIM_Command(32'd94346400);
PIM_Command(32'd75665057);
PIM_Command(32'd75534498);
PIM_Command(32'd94544291);
PIM_Command(32'd75730340);
PIM_Command(32'd94675365);
PIM_Command(32'd93948838);
PIM_Command(32'd94086567);
PIM_Command(32'd94282664);
PIM_Command(32'd94414249);
PIM_Command(32'd94806954);
PIM_Command(32'd94867883);
PIM_Command(32'd94933932);
PIM_Command(32'd94999725);
PIM_Command(32'd95071150);
PIM_Command(32'd78294191);
PIM_Command(32'd95268784);
PIM_Command(32'd78557361);
PIM_Command(32'd95529906);
PIM_Command(32'd95202739);
PIM_Command(32'd95137716);
PIM_Command(32'd78951349);
PIM_Command(32'd95792566);
PIM_Command(32'd95205047);
PIM_Command(32'd95467192);
PIM_Command(32'd78493881);
PIM_Command(32'd96057274);
PIM_Command(32'd95467963);
PIM_Command(32'd78822332);
PIM_Command(32'd95337661);
PIM_Command(32'd96320190);
PIM_Command(32'd95598271);
PIM_Command(32'd95600064);
PIM_Command(32'd95861441);
PIM_Command(32'd96452290);
PIM_Command(32'd79792835);
PIM_Command(32'd79334596);
PIM_Command(32'd79063237);
PIM_Command(32'd79729350);
PIM_Command(32'd79529159);
PIM_Command(32'd78811080);
PIM_Command(32'd79662793);
PIM_Command(32'd79859914);
PIM_Command(32'd79597003);
PIM_Command(32'd79791820);
PIM_Command(32'd79333837);
PIM_Command(32'd79070670);
PIM_Command(32'd79725007);
PIM_Command(32'd79530192);
PIM_Command(32'd78809041);
PIM_Command(32'd79659730);
PIM_Command(32'd79855827);
PIM_Command(32'd79594452);
PIM_Command(32'd97702869);
PIM_Command(32'd97375702);
PIM_Command(32'd97310423);
PIM_Command(32'd96716248);
PIM_Command(32'd96781273);
PIM_Command(32'd96913370);
PIM_Command(32'd97507547);
PIM_Command(32'd97180380);
PIM_Command(32'd97246173);
PIM_Command(32'd98360798);
PIM_Command(32'd98228703);
PIM_Command(32'd96913632);
PIM_Command(32'd97572321);
PIM_Command(32'd98099426);
PIM_Command(32'd98033516);
PIM_Command(32'd97115363);
PIM_Command(32'd97640164);
PIM_Command(32'd98689765);
PIM_Command(32'd298837352);
PIM_Command(32'd97706982);
PIM_Command(32'd97963751);
PIM_Command(32'd98034543);
PIM_Command(32'd299820393);
PIM_Command(32'd98724971);
PIM_Command(32'd292348782);
PIM_Command(32'd98887400);
PIM_Command(32'd300471405);
PIM_Command(32'd99083370);
PIM_Command(32'd91517568);
PIM_Command(32'd91713921);
PIM_Command(32'd91714690);
PIM_Command(32'd91714179);
PIM_Command(32'd91649429);
PIM_Command(32'd93679748);
PIM_Command(32'd92566661);
PIM_Command(32'd92373126);
PIM_Command(32'd92567431);
PIM_Command(32'd92565896);
PIM_Command(32'd92832649);
PIM_Command(32'd91457174);
PIM_Command(32'd93745802);
PIM_Command(32'd93746827);
PIM_Command(32'd92958860);
PIM_Command(32'd92968333);
PIM_Command(32'd93029006);
PIM_Command(32'd91262607);
PIM_Command(32'd93163152);
PIM_Command(32'd93160337);
PIM_Command(32'd93687442);
PIM_Command(32'd92377747);
PIM_Command(32'd91722388);
PIM_Command(32'd75926167);
PIM_Command(32'd76123288);
PIM_Command(32'd93886361);
PIM_Command(32'd75853978);
PIM_Command(32'd94017435);
PIM_Command(32'd75600540);
PIM_Command(32'd76055709);
PIM_Command(32'd94215326);
PIM_Command(32'd75992991);
PIM_Command(32'd94346400);
PIM_Command(32'd75665057);
PIM_Command(32'd75534498);
PIM_Command(32'd94544291);
PIM_Command(32'd75730340);
PIM_Command(32'd94675365);
PIM_Command(32'd93948838);
PIM_Command(32'd94086567);
PIM_Command(32'd94282664);
PIM_Command(32'd94414249);
PIM_Command(32'd94806954);
PIM_Command(32'd94867883);
PIM_Command(32'd94933932);
PIM_Command(32'd94999725);
PIM_Command(32'd95071150);
PIM_Command(32'd78294191);
PIM_Command(32'd95268784);
PIM_Command(32'd78557361);
PIM_Command(32'd95529906);
PIM_Command(32'd95202739);
PIM_Command(32'd95137716);
PIM_Command(32'd78951349);
PIM_Command(32'd95792566);
PIM_Command(32'd95205047);
PIM_Command(32'd95467192);
PIM_Command(32'd78493881);
PIM_Command(32'd96057274);
PIM_Command(32'd95467963);
PIM_Command(32'd78822332);
PIM_Command(32'd95337661);
PIM_Command(32'd96320190);
PIM_Command(32'd95598271);
PIM_Command(32'd95600064);
PIM_Command(32'd95861441);
PIM_Command(32'd96452290);
PIM_Command(32'd79792835);
PIM_Command(32'd79334596);
PIM_Command(32'd79065285);
PIM_Command(32'd79729350);
PIM_Command(32'd79529159);
PIM_Command(32'd78811080);
PIM_Command(32'd79662793);
PIM_Command(32'd79859914);
PIM_Command(32'd79597003);
PIM_Command(32'd79791820);
PIM_Command(32'd79333837);
PIM_Command(32'd79070670);
PIM_Command(32'd79725007);
PIM_Command(32'd79530192);
PIM_Command(32'd78809041);
PIM_Command(32'd79659730);
PIM_Command(32'd79855827);
PIM_Command(32'd79594452);
PIM_Command(32'd97702869);
PIM_Command(32'd97375702);
PIM_Command(32'd97310423);
PIM_Command(32'd96716248);
PIM_Command(32'd96781273);
PIM_Command(32'd96913370);
PIM_Command(32'd97507547);
PIM_Command(32'd97180380);
PIM_Command(32'd97246173);
PIM_Command(32'd98360798);
PIM_Command(32'd98228703);
PIM_Command(32'd96913632);
PIM_Command(32'd97572321);
PIM_Command(32'd98099426);
PIM_Command(32'd98033524);
PIM_Command(32'd97115363);
PIM_Command(32'd97640164);
PIM_Command(32'd98689765);
PIM_Command(32'd298837360);
PIM_Command(32'd97706982);
PIM_Command(32'd97963751);
PIM_Command(32'd98034551);
PIM_Command(32'd299820401);
PIM_Command(32'd98727027);
PIM_Command(32'd292873078);
PIM_Command(32'd98887400);
PIM_Command(32'd300471413);
PIM_Command(32'd99083378);
PIM_Command(32'd92043904);
PIM_Command(32'd92240257);
PIM_Command(32'd92241026);
PIM_Command(32'd92240515);
PIM_Command(32'd92175765);
PIM_Command(32'd93681796);
PIM_Command(32'd92568709);
PIM_Command(32'd92373126);
PIM_Command(32'd92569479);
PIM_Command(32'd92567944);
PIM_Command(32'd92832649);
PIM_Command(32'd91981462);
PIM_Command(32'd93747850);
PIM_Command(32'd93748875);
PIM_Command(32'd92960908);
PIM_Command(32'd92968333);
PIM_Command(32'd93029006);
PIM_Command(32'd91786895);
PIM_Command(32'd93163152);
PIM_Command(32'd93160337);
PIM_Command(32'd93687442);
PIM_Command(32'd92377747);
PIM_Command(32'd92246676);
PIM_Command(32'd75926167);
PIM_Command(32'd76123288);
PIM_Command(32'd93886361);
PIM_Command(32'd75856026);
PIM_Command(32'd94017435);
PIM_Command(32'd75600540);
PIM_Command(32'd76055709);
PIM_Command(32'd94215326);
PIM_Command(32'd75992991);
PIM_Command(32'd94346400);
PIM_Command(32'd75665057);
PIM_Command(32'd75534498);
PIM_Command(32'd94544291);
PIM_Command(32'd75730340);
PIM_Command(32'd94675365);
PIM_Command(32'd93948838);
PIM_Command(32'd94086567);
PIM_Command(32'd94282664);
PIM_Command(32'd94414249);
PIM_Command(32'd94806954);
PIM_Command(32'd94867883);
PIM_Command(32'd94933932);
PIM_Command(32'd94999725);
PIM_Command(32'd95071150);
PIM_Command(32'd78294191);
PIM_Command(32'd95268784);
PIM_Command(32'd78557361);
PIM_Command(32'd95529906);
PIM_Command(32'd95202739);
PIM_Command(32'd95137716);
PIM_Command(32'd78951349);
PIM_Command(32'd95792566);
PIM_Command(32'd95205047);
PIM_Command(32'd95467192);
PIM_Command(32'd78493881);
PIM_Command(32'd96057274);
PIM_Command(32'd95467963);
PIM_Command(32'd78822332);
PIM_Command(32'd95337661);
PIM_Command(32'd96320190);
PIM_Command(32'd95598271);
PIM_Command(32'd95600064);
PIM_Command(32'd95861441);
PIM_Command(32'd96452290);
PIM_Command(32'd79792835);
PIM_Command(32'd79334596);
PIM_Command(32'd79067333);
PIM_Command(32'd79729350);
PIM_Command(32'd79529159);
PIM_Command(32'd78811080);
PIM_Command(32'd79662793);
PIM_Command(32'd79859914);
PIM_Command(32'd79597003);
PIM_Command(32'd79791820);
PIM_Command(32'd79333837);
PIM_Command(32'd79070670);
PIM_Command(32'd79725007);
PIM_Command(32'd79530192);
PIM_Command(32'd78809041);
PIM_Command(32'd79659730);
PIM_Command(32'd79855827);
PIM_Command(32'd79594452);
PIM_Command(32'd97702869);
PIM_Command(32'd97375702);
PIM_Command(32'd97310423);
PIM_Command(32'd96716248);
PIM_Command(32'd96781273);
PIM_Command(32'd96913370);
PIM_Command(32'd97507547);
PIM_Command(32'd97180380);
PIM_Command(32'd97246173);
PIM_Command(32'd98360798);
PIM_Command(32'd98228703);
PIM_Command(32'd96913632);
PIM_Command(32'd97572321);
PIM_Command(32'd98099426);
PIM_Command(32'd98033532);
PIM_Command(32'd97115363);
PIM_Command(32'd97640164);
PIM_Command(32'd98689765);
PIM_Command(32'd298837368);
PIM_Command(32'd97706982);
PIM_Command(32'd97963751);
PIM_Command(32'd98034559);
PIM_Command(32'd299820409);
PIM_Command(32'd98729083);
PIM_Command(32'd293397374);
PIM_Command(32'd98887400);
PIM_Command(32'd300471421);
PIM_Command(32'd99083386);


endtask



task MC();


PIM_Command(32'd83896480);
PIM_Command(32'd89159841);
PIM_Command(32'd83962274);
PIM_Command(32'd89225635);
PIM_Command(32'd84028068);
PIM_Command(32'd89291429);
PIM_Command(32'd84093862);
PIM_Command(32'd89357223);
PIM_Command(32'd84159656);
PIM_Command(32'd89423017);
PIM_Command(32'd84225450);
PIM_Command(32'd89488811);
PIM_Command(32'd84291244);
PIM_Command(32'd89554605);
PIM_Command(32'd89620398);
PIM_Command(32'd84357039);
PIM_Command(32'd86548912);
PIM_Command(32'd95400064);
PIM_Command(32'd84367281);
PIM_Command(32'd91791538);
PIM_Command(32'd95335056);
PIM_Command(32'd94474419);
PIM_Command(32'd95531928);
PIM_Command(32'd91991732);
PIM_Command(32'd94404789);
PIM_Command(32'd95532424);
PIM_Command(32'd94745782);
PIM_Command(32'd94811795);
PIM_Command(32'd86749111);
PIM_Command(32'd94877624);
PIM_Command(32'd94681219);
PIM_Command(32'd84038329);
PIM_Command(32'd95533498);
PIM_Command(32'd95008699);
PIM_Command(32'd94942396);
PIM_Command(32'd86680253);
PIM_Command(32'd94748034);
PIM_Command(32'd91923390);
PIM_Command(32'd94682770);
PIM_Command(32'd86604223);
PIM_Command(32'd96059328);
PIM_Command(32'd96387210);
PIM_Command(32'd96321690);
PIM_Command(32'd83997377);
PIM_Command(32'd92187586);
PIM_Command(32'd95208086);
PIM_Command(32'd86945219);
PIM_Command(32'd95077254);
PIM_Command(32'd84235716);
PIM_Command(32'd92189125);
PIM_Command(32'd89239750);
PIM_Command(32'd86878407);
PIM_Command(32'd95143813);
PIM_Command(32'd86820040);
PIM_Command(32'd92121545);
PIM_Command(32'd95078805);
PIM_Command(32'd92063946);
PIM_Command(32'd97110669);
PIM_Command(32'd96979613);
PIM_Command(32'd87010507);
PIM_Command(32'd95341447);
PIM_Command(32'd86951372);
PIM_Command(32'd97242271);
PIM_Command(32'd92253645);
PIM_Command(32'd97308047);
PIM_Command(32'd95407511);
PIM_Command(32'd95208654);
PIM_Command(32'd92720782);
PIM_Command(32'd96453071);
PIM_Command(32'd95670161);
PIM_Command(32'd94798800);
PIM_Command(32'd96129163);
PIM_Command(32'd94553809);
PIM_Command(32'd93901209);
PIM_Command(32'd94868434);
PIM_Command(32'd96129691);
PIM_Command(32'd89575123);
PIM_Command(32'd95146910);
PIM_Command(32'd89373908);
PIM_Command(32'd92066964);
PIM_Command(32'd84130773);
PIM_Command(32'd86824324);
PIM_Command(32'd94618070);
PIM_Command(32'd92853897);
PIM_Command(32'd95797207);
PIM_Command(32'd96917377);
PIM_Command(32'd84193752);
PIM_Command(32'd89381081);
PIM_Command(32'd96197004);
PIM_Command(32'd84131034);
PIM_Command(32'd95541979);
PIM_Command(32'd89447324);
PIM_Command(32'd86001856);
PIM_Command(32'd91232449);
PIM_Command(32'd86067650);
PIM_Command(32'd91298243);
PIM_Command(32'd86133444);
PIM_Command(32'd91364037);
PIM_Command(32'd86199238);
PIM_Command(32'd91429831);
PIM_Command(32'd86265032);
PIM_Command(32'd91495625);
PIM_Command(32'd86330826);
PIM_Command(32'd91561419);
PIM_Command(32'd86396620);
PIM_Command(32'd91627213);
PIM_Command(32'd91693006);
PIM_Command(32'd86462415);
PIM_Command(32'd88654288);
PIM_Command(32'd97505440);
PIM_Command(32'd86472657);
PIM_Command(32'd85508306);
PIM_Command(32'd97440432);
PIM_Command(32'd96579795);
PIM_Command(32'd97637304);
PIM_Command(32'd85708500);
PIM_Command(32'd96510165);
PIM_Command(32'd97637800);
PIM_Command(32'd96851158);
PIM_Command(32'd96917171);
PIM_Command(32'd88854487);
PIM_Command(32'd96983000);
PIM_Command(32'd96786595);
PIM_Command(32'd86143705);
PIM_Command(32'd97638874);
PIM_Command(32'd97114075);
PIM_Command(32'd97047772);
PIM_Command(32'd88785629);
PIM_Command(32'd96853410);
PIM_Command(32'd85640158);
PIM_Command(32'd96788146);
PIM_Command(32'd88676831);
PIM_Command(32'd98164704);
PIM_Command(32'd98492586);
PIM_Command(32'd98427066);
PIM_Command(32'd86102753);
PIM_Command(32'd85904354);
PIM_Command(32'd97313462);
PIM_Command(32'd89050595);
PIM_Command(32'd97182630);
PIM_Command(32'd86341092);
PIM_Command(32'd85905893);
PIM_Command(32'd91345126);
PIM_Command(32'd88983783);
PIM_Command(32'd97249189);
PIM_Command(32'd88925416);
PIM_Command(32'd85838313);
PIM_Command(32'd97184181);
PIM_Command(32'd85780714);
PIM_Command(32'd99216045);
PIM_Command(32'd99084989);
PIM_Command(32'd89115883);
PIM_Command(32'd97446823);
PIM_Command(32'd89056748);
PIM_Command(32'd99347647);
PIM_Command(32'd85970413);
PIM_Command(32'd99413423);
PIM_Command(32'd97512887);
PIM_Command(32'd97314030);
PIM_Command(32'd94826158);
PIM_Command(32'd98558447);
PIM_Command(32'd97775537);
PIM_Command(32'd96904176);
PIM_Command(32'd98234539);
PIM_Command(32'd96659185);
PIM_Command(32'd96006585);
PIM_Command(32'd96973810);
PIM_Command(32'd98235067);
PIM_Command(32'd91680499);
PIM_Command(32'd97252286);
PIM_Command(32'd91479284);
PIM_Command(32'd85783732);
PIM_Command(32'd86236149);
PIM_Command(32'd88929700);
PIM_Command(32'd96723446);
PIM_Command(32'd94959273);
PIM_Command(32'd97902583);
PIM_Command(32'd99022753);
PIM_Command(32'd86299128);
PIM_Command(32'd91486457);
PIM_Command(32'd98302380);
PIM_Command(32'd86236410);
PIM_Command(32'd97647355);
PIM_Command(32'd91552700);
PIM_Command(32'd88107232);
PIM_Command(32'd84949217);
PIM_Command(32'd88173026);
PIM_Command(32'd85015011);
PIM_Command(32'd88238820);
PIM_Command(32'd85080805);
PIM_Command(32'd88304614);
PIM_Command(32'd85146599);
PIM_Command(32'd88370408);
PIM_Command(32'd85212393);
PIM_Command(32'd88436202);
PIM_Command(32'd85278187);
PIM_Command(32'd88501996);
PIM_Command(32'd85343981);
PIM_Command(32'd85409774);
PIM_Command(32'd88567791);
PIM_Command(32'd90759664);
PIM_Command(32'd99610816);
PIM_Command(32'd88545265);
PIM_Command(32'd87613682);
PIM_Command(32'd99545808);
PIM_Command(32'd98685171);
PIM_Command(32'd99742680);
PIM_Command(32'd87813876);
PIM_Command(32'd98615541);
PIM_Command(32'd99743176);
PIM_Command(32'd98956534);
PIM_Command(32'd99022547);
PIM_Command(32'd90959863);
PIM_Command(32'd99088376);
PIM_Command(32'd98891971);
PIM_Command(32'd88216313);
PIM_Command(32'd99744250);
PIM_Command(32'd99219451);
PIM_Command(32'd99153148);
PIM_Command(32'd90891005);
PIM_Command(32'd98958786);
PIM_Command(32'd87745534);
PIM_Command(32'd98893522);
PIM_Command(32'd90782207);
PIM_Command(32'd100269824);
PIM_Command(32'd100532426);
PIM_Command(32'd100466906);
PIM_Command(32'd88207873);
PIM_Command(32'd88009474);
PIM_Command(32'd99353302);
PIM_Command(32'd91155715);
PIM_Command(32'd99222470);
PIM_Command(32'd88413444);
PIM_Command(32'd88011013);
PIM_Command(32'd85061638);
PIM_Command(32'd91088903);
PIM_Command(32'd99289029);
PIM_Command(32'd90965032);
PIM_Command(32'd87943465);
PIM_Command(32'd99232213);
PIM_Command(32'd87828522);
PIM_Command(32'd86584013);
PIM_Command(32'd84355805);
PIM_Command(32'd91221035);
PIM_Command(32'd99494855);
PIM_Command(32'd91096364);
PIM_Command(32'd86715615);
PIM_Command(32'd88075565);
PIM_Command(32'd86781391);
PIM_Command(32'd99560919);
PIM_Command(32'd99353646);
PIM_Command(32'd96874190);
PIM_Command(32'd100598063);
PIM_Command(32'd99823569);
PIM_Command(32'd99009360);
PIM_Command(32'd100290763);
PIM_Command(32'd98698833);
PIM_Command(32'd98062809);
PIM_Command(32'd99078994);
PIM_Command(32'd100291291);
PIM_Command(32'd85339731);
PIM_Command(32'd99308510);
PIM_Command(32'd85195860);
PIM_Command(32'd87839956);
PIM_Command(32'd88341333);
PIM_Command(32'd90985924);
PIM_Command(32'd98763094);
PIM_Command(32'd97015497);
PIM_Command(32'd100007767);
PIM_Command(32'd84301761);
PIM_Command(32'd88404344);
PIM_Command(32'd85162105);
PIM_Command(32'd100366796);
PIM_Command(32'd88341626);
PIM_Command(32'd99711611);
PIM_Command(32'd85228508);
PIM_Command(32'd90179584);
PIM_Command(32'd87054337);
PIM_Command(32'd90245378);
PIM_Command(32'd87120131);
PIM_Command(32'd90311172);
PIM_Command(32'd87185925);
PIM_Command(32'd90376966);
PIM_Command(32'd87251719);
PIM_Command(32'd90442792);
PIM_Command(32'd87317545);
PIM_Command(32'd90508586);
PIM_Command(32'd87383339);
PIM_Command(32'd90574380);
PIM_Command(32'd87449133);
PIM_Command(32'd87514926);
PIM_Command(32'd90640175);
PIM_Command(32'd84410704);
PIM_Command(32'd86986976);
PIM_Command(32'd90650449);
PIM_Command(32'd89653330);
PIM_Command(32'd86921968);
PIM_Command(32'd84013139);
PIM_Command(32'd89215992);
PIM_Command(32'd89861716);
PIM_Command(32'd83943509);
PIM_Command(32'd89216488);
PIM_Command(32'd84235350);
PIM_Command(32'd84301555);
PIM_Command(32'd84619095);
PIM_Command(32'd84367224);
PIM_Command(32'd84179171);
PIM_Command(32'd90321529);
PIM_Command(32'd89225594);
PIM_Command(32'd86595451);
PIM_Command(32'd86529148);
PIM_Command(32'd84542077);
PIM_Command(32'd84245986);
PIM_Command(32'd89785214);
PIM_Command(32'd84180722);
PIM_Command(32'd84498815);
PIM_Command(32'd91848480);
PIM_Command(32'd92152042);
PIM_Command(32'd92086522);
PIM_Command(32'd90264097);
PIM_Command(32'd90057506);
PIM_Command(32'd86778614);
PIM_Command(32'd84815139);
PIM_Command(32'd86647782);
PIM_Command(32'd90518820);
PIM_Command(32'd90067237);
PIM_Command(32'd87117862);
PIM_Command(32'd84748327);
PIM_Command(32'd86714341);
PIM_Command(32'd84681800);
PIM_Command(32'd89991497);
PIM_Command(32'd86657525);
PIM_Command(32'd89933898);
PIM_Command(32'd88689389);
PIM_Command(32'd86461181);
PIM_Command(32'd84880459);
PIM_Command(32'd86920167);
PIM_Command(32'd84813132);
PIM_Command(32'd88820991);
PIM_Command(32'd90123597);
PIM_Command(32'd88886767);
PIM_Command(32'd86986231);
PIM_Command(32'd86778958);
PIM_Command(32'd98979566);
PIM_Command(32'd92217679);
PIM_Command(32'd89346033);
PIM_Command(32'd84337520);
PIM_Command(32'd91910379);
PIM_Command(32'd84026993);
PIM_Command(32'd100168185);
PIM_Command(32'd84407154);
PIM_Command(32'd91910907);
PIM_Command(32'd87445107);
PIM_Command(32'd86733822);
PIM_Command(32'd87260276);
PIM_Command(32'd89945332);
PIM_Command(32'd90405749);
PIM_Command(32'd84702692);
PIM_Command(32'd84091254);
PIM_Command(32'd99120873);
PIM_Command(32'd89489271);
PIM_Command(32'd86407137);
PIM_Command(32'd90460440);
PIM_Command(32'd87234585);
PIM_Command(32'd91953644);
PIM_Command(32'd90405914);
PIM_Command(32'd89201179);
PIM_Command(32'd87301116);



endtask

task inv_MC();

PIM_Command(32'd83888264);
PIM_Command(32'd84940937);
PIM_Command(32'd83954058);
PIM_Command(32'd85006731);
PIM_Command(32'd84019852);
PIM_Command(32'd85072525);
PIM_Command(32'd84085646);
PIM_Command(32'd85138319);
PIM_Command(32'd84151440);
PIM_Command(32'd85204113);
PIM_Command(32'd84217234);
PIM_Command(32'd85269907);
PIM_Command(32'd84283028);
PIM_Command(32'd85335701);
PIM_Command(32'd85401494);
PIM_Command(32'd84348823);
PIM_Command(32'd84445592);
PIM_Command(32'd93821056);
PIM_Command(32'd84350873);
PIM_Command(32'd85493914);
PIM_Command(32'd93756112);
PIM_Command(32'd92917915);
PIM_Command(32'd93953016);
PIM_Command(32'd85694108);
PIM_Command(32'd92831901);
PIM_Command(32'd93953448);
PIM_Command(32'd93166750);
PIM_Command(32'd93232851);
PIM_Command(32'd84645791);
PIM_Command(32'd93298592);
PIM_Command(32'd93102211);
PIM_Command(32'd84021921);
PIM_Command(32'd93954466);
PIM_Command(32'd93429667);
PIM_Command(32'd93363364);
PIM_Command(32'd84576933);
PIM_Command(32'd93169026);
PIM_Command(32'd85625766);
PIM_Command(32'd93103826);
PIM_Command(32'd84482471);
PIM_Command(32'd94480304);
PIM_Command(32'd94810282);
PIM_Command(32'd94744826);
PIM_Command(32'd83991217);
PIM_Command(32'd85889970);
PIM_Command(32'd93631190);
PIM_Command(32'd84841907);
PIM_Command(32'd93500294);
PIM_Command(32'd84219316);
PIM_Command(32'd85891509);
PIM_Command(32'd85039286);
PIM_Command(32'd84775095);
PIM_Command(32'd93566853);
PIM_Command(32'd84718776);
PIM_Command(32'd85823929);
PIM_Command(32'd93501909);
PIM_Command(32'd85768378);
PIM_Command(32'd96058029);
PIM_Command(32'd95927037);
PIM_Command(32'd84907195);
PIM_Command(32'd93764487);
PIM_Command(32'd84850108);
PIM_Command(32'd96189695);
PIM_Command(32'd85956029);
PIM_Command(32'd96255407);
PIM_Command(32'd93830615);
PIM_Command(32'd93631678);
PIM_Command(32'd92716718);
PIM_Command(32'd94876095);
PIM_Command(32'd94093265);
PIM_Command(32'd93225920);
PIM_Command(32'd94552235);
PIM_Command(32'd92976833);
PIM_Command(32'd100188665);
PIM_Command(32'd93311938);
PIM_Command(32'd94552827);
PIM_Command(32'd85376707);
PIM_Command(32'd93570046);
PIM_Command(32'd85173444);
PIM_Command(32'd85771476);
PIM_Command(32'd84124613);
PIM_Command(32'd84723076);
PIM_Command(32'd93041094);
PIM_Command(32'd94946985);
PIM_Command(32'd94218183);
PIM_Command(32'd95864705);
PIM_Command(32'd84187592);
PIM_Command(32'd85182665);
PIM_Command(32'd94620076);
PIM_Command(32'd84124874);
PIM_Command(32'd93965003);
PIM_Command(32'd85249020);
PIM_Command(32'd92317832);
PIM_Command(32'd97581193);
PIM_Command(32'd92383626);
PIM_Command(32'd97646987);
PIM_Command(32'd92449420);
PIM_Command(32'd97712781);
PIM_Command(32'd92515214);
PIM_Command(32'd97778575);
PIM_Command(32'd92581008);
PIM_Command(32'd97844369);
PIM_Command(32'd92646802);
PIM_Command(32'd97910163);
PIM_Command(32'd92712596);
PIM_Command(32'd97975957);
PIM_Command(32'd98041750);
PIM_Command(32'd92778391);
PIM_Command(32'd94931352);
PIM_Command(32'd93820928);
PIM_Command(32'd92788633);
PIM_Command(32'd100173978);
PIM_Command(32'd93755920);
PIM_Command(32'd92868763);
PIM_Command(32'd93952792);
PIM_Command(32'd100374172);
PIM_Command(32'd92799133);
PIM_Command(32'd93953288);
PIM_Command(32'd93166750);
PIM_Command(32'd93232659);
PIM_Command(32'd95131551);
PIM_Command(32'd93298592);
PIM_Command(32'd93102083);
PIM_Command(32'd92459681);
PIM_Command(32'd93954466);
PIM_Command(32'd93429667);
PIM_Command(32'd93363364);
PIM_Command(32'd95062693);
PIM_Command(32'd93168898);
PIM_Command(32'd100305830);
PIM_Command(32'd93103634);
PIM_Command(32'd95025575);
PIM_Command(32'd94480304);
PIM_Command(32'd94810122);
PIM_Command(32'd94744602);
PIM_Command(32'd92379825);
PIM_Command(32'd100570034);
PIM_Command(32'd93630998);
PIM_Command(32'd95327667);
PIM_Command(32'd93500166);
PIM_Command(32'd92657076);
PIM_Command(32'd100571573);
PIM_Command(32'd97622198);
PIM_Command(32'd95260855);
PIM_Command(32'd93566725);
PIM_Command(32'd95204536);
PIM_Command(32'd100503993);
PIM_Command(32'd93501717);
PIM_Command(32'd100448442);
PIM_Command(32'd96057869);
PIM_Command(32'd95926813);
PIM_Command(32'd95392955);
PIM_Command(32'd93764359);
PIM_Command(32'd95335868);
PIM_Command(32'd96189471);
PIM_Command(32'd100636093);
PIM_Command(32'd96255247);
PIM_Command(32'd93830423);
PIM_Command(32'd93631678);
PIM_Command(32'd84327950);
PIM_Command(32'd94876095);
PIM_Command(32'd94093073);
PIM_Command(32'd93193152);
PIM_Command(32'd94552075);
PIM_Command(32'd92976833);
PIM_Command(32'd85508377);
PIM_Command(32'd93262786);
PIM_Command(32'd94552603);
PIM_Command(32'd97959619);
PIM_Command(32'd93569822);
PIM_Command(32'd97756356);
PIM_Command(32'd100451348);
PIM_Command(32'd92513221);
PIM_Command(32'd95208708);
PIM_Command(32'd93041094);
PIM_Command(32'd84461065);
PIM_Command(32'd94218183);
PIM_Command(32'd95864577);
PIM_Command(32'd92576200);
PIM_Command(32'd97765577);
PIM_Command(32'd94619916);
PIM_Command(32'd92513482);
PIM_Command(32'd93965003);
PIM_Command(32'd97831708);
PIM_Command(32'd83888264);
PIM_Command(32'd84940937);
PIM_Command(32'd83954058);
PIM_Command(32'd85006731);
PIM_Command(32'd84019852);
PIM_Command(32'd85072525);
PIM_Command(32'd84085646);
PIM_Command(32'd85138319);
PIM_Command(32'd84151440);
PIM_Command(32'd85204113);
PIM_Command(32'd84217234);
PIM_Command(32'd85269907);
PIM_Command(32'd84283028);
PIM_Command(32'd85335701);
PIM_Command(32'd85401494);
PIM_Command(32'd84348823);
PIM_Command(32'd84445592);
PIM_Command(32'd93821056);
PIM_Command(32'd84350873);
PIM_Command(32'd85493914);
PIM_Command(32'd93756112);
PIM_Command(32'd92917915);
PIM_Command(32'd93953016);
PIM_Command(32'd85694108);
PIM_Command(32'd92831901);
PIM_Command(32'd93953448);
PIM_Command(32'd93166750);
PIM_Command(32'd93232851);
PIM_Command(32'd84645791);
PIM_Command(32'd93298592);
PIM_Command(32'd93102211);
PIM_Command(32'd84021921);
PIM_Command(32'd93954466);
PIM_Command(32'd93429667);
PIM_Command(32'd93363364);
PIM_Command(32'd84576933);
PIM_Command(32'd93169026);
PIM_Command(32'd85625766);
PIM_Command(32'd93103826);
PIM_Command(32'd84482471);
PIM_Command(32'd94480304);
PIM_Command(32'd94810282);
PIM_Command(32'd94744826);
PIM_Command(32'd83991217);
PIM_Command(32'd85889970);
PIM_Command(32'd93631190);
PIM_Command(32'd84841907);
PIM_Command(32'd93500294);
PIM_Command(32'd84219316);
PIM_Command(32'd85891509);
PIM_Command(32'd85039286);
PIM_Command(32'd84775095);
PIM_Command(32'd93566853);
PIM_Command(32'd84718776);
PIM_Command(32'd85823929);
PIM_Command(32'd93501909);
PIM_Command(32'd85768378);
PIM_Command(32'd96058029);
PIM_Command(32'd95927037);
PIM_Command(32'd84907195);
PIM_Command(32'd93764487);
PIM_Command(32'd84850108);
PIM_Command(32'd96189695);
PIM_Command(32'd85956029);
PIM_Command(32'd96255407);
PIM_Command(32'd93830615);
PIM_Command(32'd93631678);
PIM_Command(32'd92716718);
PIM_Command(32'd94876095);
PIM_Command(32'd94093265);
PIM_Command(32'd93225920);
PIM_Command(32'd94552235);
PIM_Command(32'd92976833);
PIM_Command(32'd100188665);
PIM_Command(32'd93311938);
PIM_Command(32'd94552827);
PIM_Command(32'd85376707);
PIM_Command(32'd93570046);
PIM_Command(32'd85173444);
PIM_Command(32'd85771476);
PIM_Command(32'd84124613);
PIM_Command(32'd84723076);
PIM_Command(32'd93041094);
PIM_Command(32'd94946985);
PIM_Command(32'd94218183);
PIM_Command(32'd95864705);
PIM_Command(32'd84187592);
PIM_Command(32'd85182665);
PIM_Command(32'd94620076);
PIM_Command(32'd84124874);
PIM_Command(32'd93965003);
PIM_Command(32'd85249020);
PIM_Command(32'd85993608);
PIM_Command(32'd87046281);
PIM_Command(32'd86059402);
PIM_Command(32'd87112075);
PIM_Command(32'd86125196);
PIM_Command(32'd87177869);
PIM_Command(32'd86190990);
PIM_Command(32'd87243663);
PIM_Command(32'd86256784);
PIM_Command(32'd87309457);
PIM_Command(32'd86322578);
PIM_Command(32'd87375251);
PIM_Command(32'd86388372);
PIM_Command(32'd87441045);
PIM_Command(32'd87506838);
PIM_Command(32'd86454167);
PIM_Command(32'd86542768);
PIM_Command(32'd93827232);
PIM_Command(32'd86456241);
PIM_Command(32'd87591090);
PIM_Command(32'd93762288);
PIM_Command(32'd92926131);
PIM_Command(32'd95531928);
PIM_Command(32'd87791284);
PIM_Command(32'd92840117);
PIM_Command(32'd95532488);
PIM_Command(32'd93172918);
PIM_Command(32'd93239027);
PIM_Command(32'd86742967);
PIM_Command(32'd93304760);
PIM_Command(32'd93108387);
PIM_Command(32'd86127289);
PIM_Command(32'd95533498);
PIM_Command(32'd93435835);
PIM_Command(32'd93369532);
PIM_Command(32'd86674109);
PIM_Command(32'd93175202);
PIM_Command(32'd87722942);
PIM_Command(32'd93110002);
PIM_Command(32'd86587839);
PIM_Command(32'd96059328);
PIM_Command(32'd96387274);
PIM_Command(32'd96321690);
PIM_Command(32'd86094529);
PIM_Command(32'd87987138);
PIM_Command(32'd93635318);
PIM_Command(32'd86939075);
PIM_Command(32'd93504422);
PIM_Command(32'd86324676);
PIM_Command(32'd87994821);
PIM_Command(32'd87142598);
PIM_Command(32'd86872263);
PIM_Command(32'd93570981);
PIM_Command(32'd86820056);
PIM_Command(32'd87921113);
PIM_Command(32'd93510133);
PIM_Command(32'd87873754);
PIM_Command(32'd98163405);
PIM_Command(32'd96983709);
PIM_Command(32'd87004379);
PIM_Command(32'd93772711);
PIM_Command(32'd86951388);
PIM_Command(32'd98294943);
PIM_Command(32'd88053213);
PIM_Command(32'd98360783);
PIM_Command(32'd93838839);
PIM_Command(32'd93635806);
PIM_Command(32'd94822094);
PIM_Command(32'd96453087);
PIM_Command(32'd95674353);
PIM_Command(32'd93234144);
PIM_Command(32'd96133323);
PIM_Command(32'd92980961);
PIM_Command(32'd93905305);
PIM_Command(32'd93320162);
PIM_Command(32'd96133787);
PIM_Command(32'd87482083);
PIM_Command(32'd93578142);
PIM_Command(32'd87276772);
PIM_Command(32'd87876852);
PIM_Command(32'd86227941);
PIM_Command(32'd86828452);
PIM_Command(32'd93045222);
PIM_Command(32'd97052361);
PIM_Command(32'd95797223);
PIM_Command(32'd96921505);
PIM_Command(32'd86290920);
PIM_Command(32'd87288041);
PIM_Command(32'd96201164);
PIM_Command(32'd86228202);
PIM_Command(32'd95546091);
PIM_Command(32'd87354268);
PIM_Command(32'd94423176);
PIM_Command(32'd99653769);
PIM_Command(32'd94488970);
PIM_Command(32'd99719563);
PIM_Command(32'd94554764);
PIM_Command(32'd99785357);
PIM_Command(32'd94620558);
PIM_Command(32'd99851151);
PIM_Command(32'd94686352);
PIM_Command(32'd99916945);
PIM_Command(32'd94752146);
PIM_Command(32'd99982739);
PIM_Command(32'd94817940);
PIM_Command(32'd100048533);
PIM_Command(32'd100114326);
PIM_Command(32'd94883735);
PIM_Command(32'd97028528);
PIM_Command(32'd93827104);
PIM_Command(32'd94894001);
PIM_Command(32'd93882546);
PIM_Command(32'd93762096);
PIM_Command(32'd92876979);
PIM_Command(32'd95531832);
PIM_Command(32'd94082740);
PIM_Command(32'd92807349);
PIM_Command(32'd95532328);
PIM_Command(32'd93172918);
PIM_Command(32'd93238835);
PIM_Command(32'd97228727);
PIM_Command(32'd93304760);
PIM_Command(32'd93108259);
PIM_Command(32'd94565049);
PIM_Command(32'd95533498);
PIM_Command(32'd93435835);
PIM_Command(32'd93369532);
PIM_Command(32'd97159869);
PIM_Command(32'd93175074);
PIM_Command(32'd94014398);
PIM_Command(32'd93109810);
PIM_Command(32'd97098175);
PIM_Command(32'd96059328);
PIM_Command(32'd96387114);
PIM_Command(32'd96321594);
PIM_Command(32'd94483137);
PIM_Command(32'd94278594);
PIM_Command(32'd93635126);
PIM_Command(32'd97424835);
PIM_Command(32'd93504294);
PIM_Command(32'd94762436);
PIM_Command(32'd94286277);
PIM_Command(32'd99725510);
PIM_Command(32'd97358023);
PIM_Command(32'd93570853);
PIM_Command(32'd97305816);
PIM_Command(32'd94212569);
PIM_Command(32'd93509941);
PIM_Command(32'd94165210);
PIM_Command(32'd98163245);
PIM_Command(32'd96983613);
PIM_Command(32'd97490139);
PIM_Command(32'd93772583);
PIM_Command(32'd97437148);
PIM_Command(32'd98294847);
PIM_Command(32'd94344669);
PIM_Command(32'd98360623);
PIM_Command(32'd93838647);
PIM_Command(32'd93635806);
PIM_Command(32'd86433326);
PIM_Command(32'd96453087);
PIM_Command(32'd95674161);
PIM_Command(32'd93201376);
PIM_Command(32'd96133163);
PIM_Command(32'd92980961);
PIM_Command(32'd87613753);
PIM_Command(32'd93271010);
PIM_Command(32'd96133691);
PIM_Command(32'd100064995);
PIM_Command(32'd93578046);
PIM_Command(32'd99859684);
PIM_Command(32'd94168116);
PIM_Command(32'd94616549);
PIM_Command(32'd97314084);
PIM_Command(32'd93045222);
PIM_Command(32'd86566441);
PIM_Command(32'd95797223);
PIM_Command(32'd96921377);
PIM_Command(32'd94679528);
PIM_Command(32'd99870953);
PIM_Command(32'd96201004);
PIM_Command(32'd94616810);
PIM_Command(32'd95546091);
PIM_Command(32'd99937084);
PIM_Command(32'd85993608);
PIM_Command(32'd87046281);
PIM_Command(32'd86059402);
PIM_Command(32'd87112075);
PIM_Command(32'd86125196);
PIM_Command(32'd87177869);
PIM_Command(32'd86190990);
PIM_Command(32'd87243663);
PIM_Command(32'd86256784);
PIM_Command(32'd87309457);
PIM_Command(32'd86322578);
PIM_Command(32'd87375251);
PIM_Command(32'd86388372);
PIM_Command(32'd87441045);
PIM_Command(32'd87506838);
PIM_Command(32'd86454167);
PIM_Command(32'd86542768);
PIM_Command(32'd93827232);
PIM_Command(32'd86456241);
PIM_Command(32'd87591090);
PIM_Command(32'd93762288);
PIM_Command(32'd92926131);
PIM_Command(32'd95531928);
PIM_Command(32'd87791284);
PIM_Command(32'd92840117);
PIM_Command(32'd95532488);
PIM_Command(32'd93172918);
PIM_Command(32'd93239027);
PIM_Command(32'd86742967);
PIM_Command(32'd93304760);
PIM_Command(32'd93108387);
PIM_Command(32'd86127289);
PIM_Command(32'd95533498);
PIM_Command(32'd93435835);
PIM_Command(32'd93369532);
PIM_Command(32'd86674109);
PIM_Command(32'd93175202);
PIM_Command(32'd87722942);
PIM_Command(32'd93110002);
PIM_Command(32'd86587839);
PIM_Command(32'd96059328);
PIM_Command(32'd96387274);
PIM_Command(32'd96321690);
PIM_Command(32'd86094529);
PIM_Command(32'd87987138);
PIM_Command(32'd93635318);
PIM_Command(32'd86939075);
PIM_Command(32'd93504422);
PIM_Command(32'd86324676);
PIM_Command(32'd87994821);
PIM_Command(32'd87142598);
PIM_Command(32'd86872263);
PIM_Command(32'd93570981);
PIM_Command(32'd86820056);
PIM_Command(32'd87921113);
PIM_Command(32'd93510133);
PIM_Command(32'd87873754);
PIM_Command(32'd98163405);
PIM_Command(32'd96983709);
PIM_Command(32'd87004379);
PIM_Command(32'd93772711);
PIM_Command(32'd86951388);
PIM_Command(32'd98294943);
PIM_Command(32'd88053213);
PIM_Command(32'd98360783);
PIM_Command(32'd93838839);
PIM_Command(32'd93635806);
PIM_Command(32'd94822094);
PIM_Command(32'd96453087);
PIM_Command(32'd95674353);
PIM_Command(32'd93234144);
PIM_Command(32'd96133323);
PIM_Command(32'd92980961);
PIM_Command(32'd93905305);
PIM_Command(32'd93320162);
PIM_Command(32'd96133787);
PIM_Command(32'd87482083);
PIM_Command(32'd93578142);
PIM_Command(32'd87276772);
PIM_Command(32'd87876852);
PIM_Command(32'd86227941);
PIM_Command(32'd86828452);
PIM_Command(32'd93045222);
PIM_Command(32'd97052361);
PIM_Command(32'd95797223);
PIM_Command(32'd96921505);
PIM_Command(32'd86290920);
PIM_Command(32'd87288041);
PIM_Command(32'd96201164);
PIM_Command(32'd86228202);
PIM_Command(32'd95546091);
PIM_Command(32'd87354268);
PIM_Command(32'd88098952);
PIM_Command(32'd89151625);
PIM_Command(32'd88164746);
PIM_Command(32'd89217419);
PIM_Command(32'd88230540);
PIM_Command(32'd89283213);
PIM_Command(32'd88296334);
PIM_Command(32'd89349007);
PIM_Command(32'd88362160);
PIM_Command(32'd89414833);
PIM_Command(32'd88427954);
PIM_Command(32'd89480627);
PIM_Command(32'd88493748);
PIM_Command(32'd89546421);
PIM_Command(32'd89612214);
PIM_Command(32'd88559543);
PIM_Command(32'd88639960);
PIM_Command(32'd95934656);
PIM_Command(32'd88561625);
PIM_Command(32'd89688282);
PIM_Command(32'd95869584);
PIM_Command(32'd92901595);
PIM_Command(32'd98163640);
PIM_Command(32'd89896668);
PIM_Command(32'd92848349);
PIM_Command(32'd98164200);
PIM_Command(32'd93183198);
PIM_Command(32'd93249171);
PIM_Command(32'd88848351);
PIM_Command(32'd93315040);
PIM_Command(32'd93118659);
PIM_Command(32'd88232673);
PIM_Command(32'd98165218);
PIM_Command(32'd95543267);
PIM_Command(32'd95476964);
PIM_Command(32'd88771301);
PIM_Command(32'd93185474);
PIM_Command(32'd89820134);
PIM_Command(32'd93120146);
PIM_Command(32'd88693223);
PIM_Command(32'd98690816);
PIM_Command(32'd98959594);
PIM_Command(32'd98894010);
PIM_Command(32'd88201729);
PIM_Command(32'd90092290);
PIM_Command(32'd95683222);
PIM_Command(32'd89044227);
PIM_Command(32'd95552454);
PIM_Command(32'd88429828);
PIM_Command(32'd90102021);
PIM_Command(32'd89249798);
PIM_Command(32'd88977415);
PIM_Command(32'd95619013);
PIM_Command(32'd88867848);
PIM_Command(32'd90026249);
PIM_Command(32'd95553941);
PIM_Command(32'd89917450);
PIM_Command(32'd84478701);
PIM_Command(32'd84347581);
PIM_Command(32'd89109515);
PIM_Command(32'd95816647);
PIM_Command(32'd88999180);
PIM_Command(32'd84610239);
PIM_Command(32'd90158349);
PIM_Command(32'd84676079);
PIM_Command(32'd95882647);
PIM_Command(32'd95683598);
PIM_Command(32'd96866030);
PIM_Command(32'd99025167);
PIM_Command(32'd98242449);
PIM_Command(32'd93242128);
PIM_Command(32'd98701547);
PIM_Command(32'd92931601);
PIM_Command(32'd95949241);
PIM_Command(32'd93295378);
PIM_Command(32'd98702011);
PIM_Command(32'd89525779);
PIM_Command(32'd95622078);
PIM_Command(32'd89383956);
PIM_Command(32'd89920660);
PIM_Command(32'd88335125);
PIM_Command(32'd88872388);
PIM_Command(32'd92995862);
PIM_Command(32'd99096297);
PIM_Command(32'd98428695);
PIM_Command(32'd84285377);
PIM_Command(32'd88398104);
PIM_Command(32'd89331737);
PIM_Command(32'd98769388);
PIM_Command(32'd88335386);
PIM_Command(32'd98114075);
PIM_Command(32'd89398204);
PIM_Command(32'd96528520);
PIM_Command(32'd93370505);
PIM_Command(32'd96594314);
PIM_Command(32'd93436299);
PIM_Command(32'd96660108);
PIM_Command(32'd93502093);
PIM_Command(32'd96725902);
PIM_Command(32'd93567887);
PIM_Command(32'd96791728);
PIM_Command(32'd93633713);
PIM_Command(32'd96857522);
PIM_Command(32'd93699507);
PIM_Command(32'd96923316);
PIM_Command(32'd93765301);
PIM_Command(32'd93831094);
PIM_Command(32'd96989111);
PIM_Command(32'd99125720);
PIM_Command(32'd95934528);
PIM_Command(32'd96966617);
PIM_Command(32'd95979738);
PIM_Command(32'd95869520);
PIM_Command(32'd92885211);
PIM_Command(32'd98163544);
PIM_Command(32'd96188124);
PIM_Command(32'd92815581);
PIM_Command(32'd98164040);
PIM_Command(32'd93183198);
PIM_Command(32'd93249107);
PIM_Command(32'd99334111);
PIM_Command(32'd93315040);
PIM_Command(32'd93118531);
PIM_Command(32'd96637665);
PIM_Command(32'd98165218);
PIM_Command(32'd95543267);
PIM_Command(32'd95476964);
PIM_Command(32'd99257061);
PIM_Command(32'd93185346);
PIM_Command(32'd96111590);
PIM_Command(32'd93120082);
PIM_Command(32'd99203559);
PIM_Command(32'd98690816);
PIM_Command(32'd98959434);
PIM_Command(32'd98893914);
PIM_Command(32'd96590337);
PIM_Command(32'd96383746);
PIM_Command(32'd95683158);
PIM_Command(32'd99529987);
PIM_Command(32'd95552326);
PIM_Command(32'd96834820);
PIM_Command(32'd96393477);
PIM_Command(32'd93444102);
PIM_Command(32'd99463175);
PIM_Command(32'd95618885);
PIM_Command(32'd99353608);
PIM_Command(32'd96317705);
PIM_Command(32'd95553877);
PIM_Command(32'd96208906);
PIM_Command(32'd84478541);
PIM_Command(32'd84347485);
PIM_Command(32'd99595275);
PIM_Command(32'd95816519);
PIM_Command(32'd99484940);
PIM_Command(32'd84610143);
PIM_Command(32'd96449805);
PIM_Command(32'd84675919);
PIM_Command(32'd95882583);
PIM_Command(32'd95683598);
PIM_Command(32'd88477262);
PIM_Command(32'd99025167);
PIM_Command(32'd98242385);
PIM_Command(32'd93209360);
PIM_Command(32'd98701387);
PIM_Command(32'd92931601);
PIM_Command(32'd89657689);
PIM_Command(32'd93278994);
PIM_Command(32'd98701915);
PIM_Command(32'd93720083);
PIM_Command(32'd95621982);
PIM_Command(32'd93578260);
PIM_Command(32'd96212052);
PIM_Command(32'd96723733);
PIM_Command(32'd99358020);
PIM_Command(32'd92995862);
PIM_Command(32'd88610377);
PIM_Command(32'd98428695);
PIM_Command(32'd84285249);
PIM_Command(32'd96786712);
PIM_Command(32'd93526041);
PIM_Command(32'd98769228);
PIM_Command(32'd96723994);
PIM_Command(32'd98114075);
PIM_Command(32'd93592412);
PIM_Command(32'd88098952);
PIM_Command(32'd89151625);
PIM_Command(32'd88164746);
PIM_Command(32'd89217419);
PIM_Command(32'd88230540);
PIM_Command(32'd89283213);
PIM_Command(32'd88296334);
PIM_Command(32'd89349007);
PIM_Command(32'd88362160);
PIM_Command(32'd89414833);
PIM_Command(32'd88427954);
PIM_Command(32'd89480627);
PIM_Command(32'd88493748);
PIM_Command(32'd89546421);
PIM_Command(32'd89612214);
PIM_Command(32'd88559543);
PIM_Command(32'd88639960);
PIM_Command(32'd95934656);
PIM_Command(32'd88561625);
PIM_Command(32'd89688282);
PIM_Command(32'd95869584);
PIM_Command(32'd92901595);
PIM_Command(32'd98163640);
PIM_Command(32'd89896668);
PIM_Command(32'd92848349);
PIM_Command(32'd98164200);
PIM_Command(32'd93183198);
PIM_Command(32'd93249171);
PIM_Command(32'd88848351);
PIM_Command(32'd93315040);
PIM_Command(32'd93118659);
PIM_Command(32'd88232673);
PIM_Command(32'd98165218);
PIM_Command(32'd95543267);
PIM_Command(32'd95476964);
PIM_Command(32'd88771301);
PIM_Command(32'd93185474);
PIM_Command(32'd89820134);
PIM_Command(32'd93120146);
PIM_Command(32'd88693223);
PIM_Command(32'd98690816);
PIM_Command(32'd98959594);
PIM_Command(32'd98894010);
PIM_Command(32'd88201729);
PIM_Command(32'd90092290);
PIM_Command(32'd95683222);
PIM_Command(32'd89044227);
PIM_Command(32'd95552454);
PIM_Command(32'd88429828);
PIM_Command(32'd90102021);
PIM_Command(32'd89249798);
PIM_Command(32'd88977415);
PIM_Command(32'd95619013);
PIM_Command(32'd88867848);
PIM_Command(32'd90026249);
PIM_Command(32'd95553941);
PIM_Command(32'd89917450);
PIM_Command(32'd84478701);
PIM_Command(32'd84347581);
PIM_Command(32'd89109515);
PIM_Command(32'd95816647);
PIM_Command(32'd88999180);
PIM_Command(32'd84610239);
PIM_Command(32'd90158349);
PIM_Command(32'd84676079);
PIM_Command(32'd95882647);
PIM_Command(32'd95683598);
PIM_Command(32'd96866030);
PIM_Command(32'd99025167);
PIM_Command(32'd98242449);
PIM_Command(32'd93242128);
PIM_Command(32'd98701547);
PIM_Command(32'd92931601);
PIM_Command(32'd95949241);
PIM_Command(32'd93295378);
PIM_Command(32'd98702011);
PIM_Command(32'd89525779);
PIM_Command(32'd95622078);
PIM_Command(32'd89383956);
PIM_Command(32'd89920660);
PIM_Command(32'd88335125);
PIM_Command(32'd88872388);
PIM_Command(32'd92995862);
PIM_Command(32'd99096297);
PIM_Command(32'd98428695);
PIM_Command(32'd84285377);
PIM_Command(32'd88398104);
PIM_Command(32'd89331737);
PIM_Command(32'd98769388);
PIM_Command(32'd88335386);
PIM_Command(32'd98114075);
PIM_Command(32'd89398204);
PIM_Command(32'd90204160);
PIM_Command(32'd91256833);
PIM_Command(32'd90269954);
PIM_Command(32'd91322627);
PIM_Command(32'd90335748);
PIM_Command(32'd91388421);
PIM_Command(32'd90401542);
PIM_Command(32'd91454215);
PIM_Command(32'd90467336);
PIM_Command(32'd91520009);
PIM_Command(32'd90533130);
PIM_Command(32'd91585803);
PIM_Command(32'd90598924);
PIM_Command(32'd91651597);
PIM_Command(32'd91717390);
PIM_Command(32'd90664719);
PIM_Command(32'd90702096);
PIM_Command(32'd84873440);
PIM_Command(32'd90666769);
PIM_Command(32'd91750418);
PIM_Command(32'd84808368);
PIM_Command(32'd83996691);
PIM_Command(32'd85005272);
PIM_Command(32'd91950612);
PIM_Command(32'd83943445);
PIM_Command(32'd85005704);
PIM_Command(32'd84218902);
PIM_Command(32'd84285107);
PIM_Command(32'd90902295);
PIM_Command(32'd84350744);
PIM_Command(32'd84154595);
PIM_Command(32'd90337817);
PIM_Command(32'd85006618);
PIM_Command(32'd84481819);
PIM_Command(32'd84415516);
PIM_Command(32'd90833437);
PIM_Command(32'd84221410);
PIM_Command(32'd91882270);
PIM_Command(32'd84156082);
PIM_Command(32'd90798367);
PIM_Command(32'd85532448);
PIM_Command(32'd85860490);
PIM_Command(32'd85795034);
PIM_Command(32'd90247713);
PIM_Command(32'd92146466);
PIM_Command(32'd84681398);
PIM_Command(32'd91098403);
PIM_Command(32'd84550630);
PIM_Command(32'd90535204);
PIM_Command(32'd92148005);
PIM_Command(32'd91295782);
PIM_Command(32'd91031591);
PIM_Command(32'd84617189);
PIM_Command(32'd90973224);
PIM_Command(32'd92080425);
PIM_Command(32'd84552117);
PIM_Command(32'd92022826);
PIM_Command(32'd86583949);
PIM_Command(32'd86452957);
PIM_Command(32'd91163691);
PIM_Command(32'd84814823);
PIM_Command(32'd91104556);
PIM_Command(32'd86715615);
PIM_Command(32'd92212525);
PIM_Command(32'd86781327);
PIM_Command(32'd84880823);
PIM_Command(32'd84681774);
PIM_Command(32'd98971278);
PIM_Command(32'd85926191);
PIM_Command(32'd85143473);
PIM_Command(32'd84337456);
PIM_Command(32'd85602443);
PIM_Command(32'd84026929);
PIM_Command(32'd98054617);
PIM_Command(32'd84390706);
PIM_Command(32'd85603035);
PIM_Command(32'd91631155);
PIM_Command(32'd84620254);
PIM_Command(32'd91429940);
PIM_Command(32'd92026036);
PIM_Command(32'd90381109);
PIM_Command(32'd90977764);
PIM_Command(32'd84091190);
PIM_Command(32'd92812937);
PIM_Command(32'd85270327);
PIM_Command(32'd86390753);
PIM_Command(32'd90444088);
PIM_Command(32'd91437113);
PIM_Command(32'd85670284);
PIM_Command(32'd90381370);
PIM_Command(32'd85015099);
PIM_Command(32'd91503580);
PIM_Command(32'd98600960);
PIM_Command(32'd95475713);
PIM_Command(32'd98666754);
PIM_Command(32'd95541507);
PIM_Command(32'd98732548);
PIM_Command(32'd95607301);
PIM_Command(32'd98798342);
PIM_Command(32'd95673095);
PIM_Command(32'd98864136);
PIM_Command(32'd95738889);
PIM_Command(32'd98929930);
PIM_Command(32'd95804683);
PIM_Command(32'd98995724);
PIM_Command(32'd95870477);
PIM_Command(32'd95936270);
PIM_Command(32'd99061519);
PIM_Command(32'd92799248);
PIM_Command(32'd84873312);
PIM_Command(32'd99071761);
PIM_Command(32'd98041874);
PIM_Command(32'd84808304);
PIM_Command(32'd83980307);
PIM_Command(32'd85005176);
PIM_Command(32'd98242068);
PIM_Command(32'd83910677);
PIM_Command(32'd85005672);
PIM_Command(32'd84218902);
PIM_Command(32'd84285043);
PIM_Command(32'd92999447);
PIM_Command(32'd84350744);
PIM_Command(32'd84154467);
PIM_Command(32'd98742809);
PIM_Command(32'd85006618);
PIM_Command(32'd84481819);
PIM_Command(32'd84415516);
PIM_Command(32'd92930589);
PIM_Command(32'd84221282);
PIM_Command(32'd98173726);
PIM_Command(32'd84156018);
PIM_Command(32'd92920095);
PIM_Command(32'd85532448);
PIM_Command(32'd85860458);
PIM_Command(32'd85794938);
PIM_Command(32'd98636321);
PIM_Command(32'd98437922);
PIM_Command(32'd84681334);
PIM_Command(32'd93195555);
PIM_Command(32'd84550502);
PIM_Command(32'd98940196);
PIM_Command(32'd98439461);
PIM_Command(32'd95490086);
PIM_Command(32'd93128743);
PIM_Command(32'd84617061);
PIM_Command(32'd93070376);
PIM_Command(32'd98371881);
PIM_Command(32'd84552053);
PIM_Command(32'd98314282);
PIM_Command(32'd86583917);
PIM_Command(32'd86452861);
PIM_Command(32'd93260843);
PIM_Command(32'd84814695);
PIM_Command(32'd93201708);
PIM_Command(32'd86715519);
PIM_Command(32'd98503981);
PIM_Command(32'd86781295);
PIM_Command(32'd84880759);
PIM_Command(32'd84681774);
PIM_Command(32'd90582638);
PIM_Command(32'd85926191);
PIM_Command(32'd85143409);
PIM_Command(32'd84304688);
PIM_Command(32'd85602411);
PIM_Command(32'd84026929);
PIM_Command(32'd91763065);
PIM_Command(32'd84374322);
PIM_Command(32'd85602939);
PIM_Command(32'd95825459);
PIM_Command(32'd84620158);
PIM_Command(32'd95624244);
PIM_Command(32'd98317428);
PIM_Command(32'd98769717);
PIM_Command(32'd93074788);
PIM_Command(32'd84091190);
PIM_Command(32'd90715753);
PIM_Command(32'd85270327);
PIM_Command(32'd86390625);
PIM_Command(32'd98832696);
PIM_Command(32'd95631417);
PIM_Command(32'd85670252);
PIM_Command(32'd98769978);
PIM_Command(32'd85015099);
PIM_Command(32'd95697788);
PIM_Command(32'd90204160);
PIM_Command(32'd91256833);
PIM_Command(32'd90269954);
PIM_Command(32'd91322627);
PIM_Command(32'd90335748);
PIM_Command(32'd91388421);
PIM_Command(32'd90401542);
PIM_Command(32'd91454215);
PIM_Command(32'd90467336);
PIM_Command(32'd91520009);
PIM_Command(32'd90533130);
PIM_Command(32'd91585803);
PIM_Command(32'd90598924);
PIM_Command(32'd91651597);
PIM_Command(32'd91717390);
PIM_Command(32'd90664719);
PIM_Command(32'd90702096);
PIM_Command(32'd84873440);
PIM_Command(32'd90666769);
PIM_Command(32'd91750418);
PIM_Command(32'd84808368);
PIM_Command(32'd83996691);
PIM_Command(32'd85005272);
PIM_Command(32'd91950612);
PIM_Command(32'd83943445);
PIM_Command(32'd85005704);
PIM_Command(32'd84218902);
PIM_Command(32'd84285107);
PIM_Command(32'd90902295);
PIM_Command(32'd84350744);
PIM_Command(32'd84154595);
PIM_Command(32'd90337817);
PIM_Command(32'd85006618);
PIM_Command(32'd84481819);
PIM_Command(32'd84415516);
PIM_Command(32'd90833437);
PIM_Command(32'd84221410);
PIM_Command(32'd91882270);
PIM_Command(32'd84156082);
PIM_Command(32'd90798367);
PIM_Command(32'd85532448);
PIM_Command(32'd85860490);
PIM_Command(32'd85795034);
PIM_Command(32'd90247713);
PIM_Command(32'd92146466);
PIM_Command(32'd84681398);
PIM_Command(32'd91098403);
PIM_Command(32'd84550630);
PIM_Command(32'd90535204);
PIM_Command(32'd92148005);
PIM_Command(32'd91295782);
PIM_Command(32'd91031591);
PIM_Command(32'd84617189);
PIM_Command(32'd90973224);
PIM_Command(32'd92080425);
PIM_Command(32'd84552117);
PIM_Command(32'd92022826);
PIM_Command(32'd86583949);
PIM_Command(32'd86452957);
PIM_Command(32'd91163691);
PIM_Command(32'd84814823);
PIM_Command(32'd91104556);
PIM_Command(32'd86715615);
PIM_Command(32'd92212525);
PIM_Command(32'd86781327);
PIM_Command(32'd84880823);
PIM_Command(32'd84681774);
PIM_Command(32'd98971278);
PIM_Command(32'd85926191);
PIM_Command(32'd85143473);
PIM_Command(32'd84337456);
PIM_Command(32'd85602443);
PIM_Command(32'd84026929);
PIM_Command(32'd98054617);
PIM_Command(32'd84390706);
PIM_Command(32'd85603035);
PIM_Command(32'd91631155);
PIM_Command(32'd84620254);
PIM_Command(32'd91429940);
PIM_Command(32'd92026036);
PIM_Command(32'd90381109);
PIM_Command(32'd90977764);
PIM_Command(32'd84091190);
PIM_Command(32'd92812937);
PIM_Command(32'd85270327);
PIM_Command(32'd86390753);
PIM_Command(32'd90444088);
PIM_Command(32'd91437113);
PIM_Command(32'd85670284);
PIM_Command(32'd90381370);
PIM_Command(32'd85015099);
PIM_Command(32'd91503580);



endtask

task inv_SBOX();

PIM_Command(32'd92767232);
PIM_Command(32'd294028289);
PIM_Command(32'd294094338);
PIM_Command(32'd92570371);
PIM_Command(32'd293830660);
PIM_Command(32'd92372997);
PIM_Command(32'd293994502);
PIM_Command(32'd83952903);
PIM_Command(32'd293602056);
PIM_Command(32'd84018185);
PIM_Command(32'd84018442);
PIM_Command(32'd84083979);
PIM_Command(32'd293929740);
PIM_Command(32'd92700941);
PIM_Command(32'd293930766);
PIM_Command(32'd84151567);
PIM_Command(32'd92472848);
PIM_Command(32'd293962257);
PIM_Command(32'd293765394);
PIM_Command(32'd293962515);
PIM_Command(32'd92737812);
PIM_Command(32'd83955989);
PIM_Command(32'd84742934);
PIM_Command(32'd84087319);
PIM_Command(32'd84481816);
PIM_Command(32'd84480537);
PIM_Command(32'd84612634);
PIM_Command(32'd67769627);
PIM_Command(32'd67110428);
PIM_Command(32'd85531421);
PIM_Command(32'd67572766);
PIM_Command(32'd85859103);
PIM_Command(32'd67835424);
PIM_Command(32'd67176481);
PIM_Command(32'd85598242);
PIM_Command(32'd68095523);
PIM_Command(32'd86188068);
PIM_Command(32'd67311653);
PIM_Command(32'd68163366);
PIM_Command(32'd86385959);
PIM_Command(32'd67242280);
PIM_Command(32'd86517033);
PIM_Command(32'd85793834);
PIM_Command(32'd85918763);
PIM_Command(32'd86122796);
PIM_Command(32'd86255917);
PIM_Command(32'd86648622);
PIM_Command(32'd86714671);
PIM_Command(32'd86779696);
PIM_Command(32'd86838321);
PIM_Command(32'd87044402);
PIM_Command(32'd70266419);
PIM_Command(32'd86979380);
PIM_Command(32'd86912821);
PIM_Command(32'd87110454);
PIM_Command(32'd70661431);
PIM_Command(32'd70529592);
PIM_Command(32'd70136121);
PIM_Command(32'd70596922);
PIM_Command(32'd87372603);
PIM_Command(32'd70201404);
PIM_Command(32'd70401085);
PIM_Command(32'd87175998);
PIM_Command(32'd86980415);
PIM_Command(32'd87702336);
PIM_Command(32'd87111745);
PIM_Command(32'd87899714);
PIM_Command(32'd88097347);
PIM_Command(32'd88031556);
PIM_Command(32'd88031301);
PIM_Command(32'd88162886);
PIM_Command(32'd88359751);
PIM_Command(32'd71701832);
PIM_Command(32'd71435849);
PIM_Command(32'd71373898);
PIM_Command(32'd71636555);
PIM_Command(32'd71305292);
PIM_Command(32'd71241293);
PIM_Command(32'd71571534);
PIM_Command(32'd71767887);
PIM_Command(32'd71502160);
PIM_Command(32'd71699025);
PIM_Command(32'd71434322);
PIM_Command(32'd71370579);
PIM_Command(32'd71633748);
PIM_Command(32'd71303509);
PIM_Command(32'd71241558);
PIM_Command(32'd71566167);
PIM_Command(32'd71766104);
PIM_Command(32'd71500377);
PIM_Command(32'd89020250);
PIM_Command(32'd89412955);
PIM_Command(32'd89151580);
PIM_Command(32'd88689757);
PIM_Command(32'd88756830);
PIM_Command(32'd88624479);
PIM_Command(32'd88823392);
PIM_Command(32'd89807713);
PIM_Command(32'd88887138);
PIM_Command(32'd89217379);
PIM_Command(32'd89349732);
PIM_Command(32'd89808229);
PIM_Command(32'd88623718);
PIM_Command(32'd88821095);
PIM_Command(32'd88823912);
PIM_Command(32'd89150825);
PIM_Command(32'd89347946);
PIM_Command(32'd89414763);
PIM_Command(32'd89743212);
PIM_Command(32'd89939309);
PIM_Command(32'd90071150);
PIM_Command(32'd89940335);
PIM_Command(32'd90268272);
PIM_Command(32'd90136945);
PIM_Command(32'd90203250);
PIM_Command(32'd90400115);
PIM_Command(32'd90467444);
PIM_Command(32'd90534517);
PIM_Command(32'd90795638);
PIM_Command(32'd90664839);
PIM_Command(32'd91453062);
PIM_Command(32'd90928517);
PIM_Command(32'd90599300);
PIM_Command(32'd91255939);
PIM_Command(32'd91058562);
PIM_Command(32'd90730625);
PIM_Command(32'd90401408);
PIM_Command(32'd93293568);
PIM_Command(32'd294554625);
PIM_Command(32'd294620674);
PIM_Command(32'd93096707);
PIM_Command(32'd294356996);
PIM_Command(32'd92899333);
PIM_Command(32'd294518790);
PIM_Command(32'd83952903);
PIM_Command(32'd294126344);
PIM_Command(32'd84018185);
PIM_Command(32'd84018442);
PIM_Command(32'd84083979);
PIM_Command(32'd294454028);
PIM_Command(32'd93227277);
PIM_Command(32'd294455054);
PIM_Command(32'd84151567);
PIM_Command(32'd92997136);
PIM_Command(32'd294488593);
PIM_Command(32'd294291730);
PIM_Command(32'd294488851);
PIM_Command(32'd93262100);
PIM_Command(32'd83955989);
PIM_Command(32'd84742934);
PIM_Command(32'd84087319);
PIM_Command(32'd84481816);
PIM_Command(32'd84480537);
PIM_Command(32'd84612634);
PIM_Command(32'd67769627);
PIM_Command(32'd67110428);
PIM_Command(32'd85531421);
PIM_Command(32'd67572766);
PIM_Command(32'd85859103);
PIM_Command(32'd67835424);
PIM_Command(32'd67176481);
PIM_Command(32'd85598242);
PIM_Command(32'd68095523);
PIM_Command(32'd86188068);
PIM_Command(32'd67311653);
PIM_Command(32'd68163366);
PIM_Command(32'd86385959);
PIM_Command(32'd67242280);
PIM_Command(32'd86517033);
PIM_Command(32'd85793834);
PIM_Command(32'd85918763);
PIM_Command(32'd86122796);
PIM_Command(32'd86255917);
PIM_Command(32'd86648622);
PIM_Command(32'd86714671);
PIM_Command(32'd86779696);
PIM_Command(32'd86838321);
PIM_Command(32'd87044402);
PIM_Command(32'd70266419);
PIM_Command(32'd86979380);
PIM_Command(32'd86912821);
PIM_Command(32'd87110454);
PIM_Command(32'd70661431);
PIM_Command(32'd70529592);
PIM_Command(32'd70136121);
PIM_Command(32'd70596922);
PIM_Command(32'd87372603);
PIM_Command(32'd70201404);
PIM_Command(32'd70401085);
PIM_Command(32'd87175998);
PIM_Command(32'd86980415);
PIM_Command(32'd87702336);
PIM_Command(32'd87111745);
PIM_Command(32'd87899714);
PIM_Command(32'd88097347);
PIM_Command(32'd88031556);
PIM_Command(32'd88031301);
PIM_Command(32'd88162886);
PIM_Command(32'd88359751);
PIM_Command(32'd71701832);
PIM_Command(32'd71435849);
PIM_Command(32'd71373898);
PIM_Command(32'd71636555);
PIM_Command(32'd71305292);
PIM_Command(32'd71241293);
PIM_Command(32'd71571534);
PIM_Command(32'd71767887);
PIM_Command(32'd71502160);
PIM_Command(32'd71699025);
PIM_Command(32'd71434322);
PIM_Command(32'd71370579);
PIM_Command(32'd71633748);
PIM_Command(32'd71303509);
PIM_Command(32'd71241558);
PIM_Command(32'd71566167);
PIM_Command(32'd71766104);
PIM_Command(32'd71500377);
PIM_Command(32'd89020250);
PIM_Command(32'd89412955);
PIM_Command(32'd89151580);
PIM_Command(32'd88689757);
PIM_Command(32'd88756830);
PIM_Command(32'd88624479);
PIM_Command(32'd88823392);
PIM_Command(32'd89807713);
PIM_Command(32'd88887138);
PIM_Command(32'd89217379);
PIM_Command(32'd89349732);
PIM_Command(32'd89808229);
PIM_Command(32'd88623718);
PIM_Command(32'd88821095);
PIM_Command(32'd88823912);
PIM_Command(32'd89150825);
PIM_Command(32'd89347946);
PIM_Command(32'd89414763);
PIM_Command(32'd89743212);
PIM_Command(32'd89939309);
PIM_Command(32'd90071150);
PIM_Command(32'd89940335);
PIM_Command(32'd90268272);
PIM_Command(32'd90136945);
PIM_Command(32'd90203250);
PIM_Command(32'd90400115);
PIM_Command(32'd90467444);
PIM_Command(32'd90534517);
PIM_Command(32'd90795638);
PIM_Command(32'd90664847);
PIM_Command(32'd91453070);
PIM_Command(32'd90928525);
PIM_Command(32'd90599308);
PIM_Command(32'd91255947);
PIM_Command(32'd91058570);
PIM_Command(32'd90730633);
PIM_Command(32'd90401416);
PIM_Command(32'd93819904);
PIM_Command(32'd295080961);
PIM_Command(32'd295147010);
PIM_Command(32'd93623043);
PIM_Command(32'd294883332);
PIM_Command(32'd93425669);
PIM_Command(32'd295043078);
PIM_Command(32'd83952903);
PIM_Command(32'd294650632);
PIM_Command(32'd84018185);
PIM_Command(32'd84018442);
PIM_Command(32'd84083979);
PIM_Command(32'd294978316);
PIM_Command(32'd93753613);
PIM_Command(32'd294979342);
PIM_Command(32'd84151567);
PIM_Command(32'd93521424);
PIM_Command(32'd295014929);
PIM_Command(32'd294818066);
PIM_Command(32'd295015187);
PIM_Command(32'd93786388);
PIM_Command(32'd83955989);
PIM_Command(32'd84742934);
PIM_Command(32'd84087319);
PIM_Command(32'd84481816);
PIM_Command(32'd84480537);
PIM_Command(32'd84612634);
PIM_Command(32'd67769627);
PIM_Command(32'd67110428);
PIM_Command(32'd85531421);
PIM_Command(32'd67572766);
PIM_Command(32'd85859103);
PIM_Command(32'd67835424);
PIM_Command(32'd67176481);
PIM_Command(32'd85598242);
PIM_Command(32'd68095523);
PIM_Command(32'd86188068);
PIM_Command(32'd67311653);
PIM_Command(32'd68163366);
PIM_Command(32'd86385959);
PIM_Command(32'd67242280);
PIM_Command(32'd86517033);
PIM_Command(32'd85793834);
PIM_Command(32'd85918763);
PIM_Command(32'd86122796);
PIM_Command(32'd86255917);
PIM_Command(32'd86648622);
PIM_Command(32'd86714671);
PIM_Command(32'd86779696);
PIM_Command(32'd86838321);
PIM_Command(32'd87044402);
PIM_Command(32'd70266419);
PIM_Command(32'd86979380);
PIM_Command(32'd86912821);
PIM_Command(32'd87110454);
PIM_Command(32'd70661431);
PIM_Command(32'd70529592);
PIM_Command(32'd70136121);
PIM_Command(32'd70596922);
PIM_Command(32'd87372603);
PIM_Command(32'd70201404);
PIM_Command(32'd70401085);
PIM_Command(32'd87175998);
PIM_Command(32'd86980415);
PIM_Command(32'd87702336);
PIM_Command(32'd87111745);
PIM_Command(32'd87899714);
PIM_Command(32'd88097347);
PIM_Command(32'd88031556);
PIM_Command(32'd88031301);
PIM_Command(32'd88162886);
PIM_Command(32'd88359751);
PIM_Command(32'd71701832);
PIM_Command(32'd71435849);
PIM_Command(32'd71373898);
PIM_Command(32'd71636555);
PIM_Command(32'd71305292);
PIM_Command(32'd71241293);
PIM_Command(32'd71571534);
PIM_Command(32'd71767887);
PIM_Command(32'd71502160);
PIM_Command(32'd71699025);
PIM_Command(32'd71434322);
PIM_Command(32'd71370579);
PIM_Command(32'd71633748);
PIM_Command(32'd71303509);
PIM_Command(32'd71241558);
PIM_Command(32'd71566167);
PIM_Command(32'd71766104);
PIM_Command(32'd71500377);
PIM_Command(32'd89020250);
PIM_Command(32'd89412955);
PIM_Command(32'd89151580);
PIM_Command(32'd88689757);
PIM_Command(32'd88756830);
PIM_Command(32'd88624479);
PIM_Command(32'd88823392);
PIM_Command(32'd89807713);
PIM_Command(32'd88887138);
PIM_Command(32'd89217379);
PIM_Command(32'd89349732);
PIM_Command(32'd89808229);
PIM_Command(32'd88623718);
PIM_Command(32'd88821095);
PIM_Command(32'd88823912);
PIM_Command(32'd89150825);
PIM_Command(32'd89347946);
PIM_Command(32'd89414763);
PIM_Command(32'd89743212);
PIM_Command(32'd89939309);
PIM_Command(32'd90071150);
PIM_Command(32'd89940335);
PIM_Command(32'd90268272);
PIM_Command(32'd90136945);
PIM_Command(32'd90203250);
PIM_Command(32'd90400115);
PIM_Command(32'd90467444);
PIM_Command(32'd90534517);
PIM_Command(32'd90795638);
PIM_Command(32'd90664855);
PIM_Command(32'd91453078);
PIM_Command(32'd90928533);
PIM_Command(32'd90599316);
PIM_Command(32'd91255955);
PIM_Command(32'd91058578);
PIM_Command(32'd90730641);
PIM_Command(32'd90401424);
PIM_Command(32'd94346240);
PIM_Command(32'd295607297);
PIM_Command(32'd295673346);
PIM_Command(32'd94149379);
PIM_Command(32'd295409668);
PIM_Command(32'd93952005);
PIM_Command(32'd295567366);
PIM_Command(32'd83952903);
PIM_Command(32'd295174920);
PIM_Command(32'd84018185);
PIM_Command(32'd84018442);
PIM_Command(32'd84083979);
PIM_Command(32'd295502604);
PIM_Command(32'd94279949);
PIM_Command(32'd295503630);
PIM_Command(32'd84151567);
PIM_Command(32'd94045712);
PIM_Command(32'd295541265);
PIM_Command(32'd295344402);
PIM_Command(32'd295541523);
PIM_Command(32'd94310676);
PIM_Command(32'd83955989);
PIM_Command(32'd84742934);
PIM_Command(32'd84087319);
PIM_Command(32'd84481816);
PIM_Command(32'd84480537);
PIM_Command(32'd84612634);
PIM_Command(32'd67769627);
PIM_Command(32'd67110428);
PIM_Command(32'd85531421);
PIM_Command(32'd67572766);
PIM_Command(32'd85859103);
PIM_Command(32'd67835424);
PIM_Command(32'd67176481);
PIM_Command(32'd85598242);
PIM_Command(32'd68095523);
PIM_Command(32'd86188068);
PIM_Command(32'd67311653);
PIM_Command(32'd68163366);
PIM_Command(32'd86385959);
PIM_Command(32'd67242280);
PIM_Command(32'd86517033);
PIM_Command(32'd85793834);
PIM_Command(32'd85918763);
PIM_Command(32'd86122796);
PIM_Command(32'd86255917);
PIM_Command(32'd86648622);
PIM_Command(32'd86714671);
PIM_Command(32'd86779696);
PIM_Command(32'd86838321);
PIM_Command(32'd87044402);
PIM_Command(32'd70266419);
PIM_Command(32'd86979380);
PIM_Command(32'd86912821);
PIM_Command(32'd87110454);
PIM_Command(32'd70661431);
PIM_Command(32'd70529592);
PIM_Command(32'd70136121);
PIM_Command(32'd70596922);
PIM_Command(32'd87372603);
PIM_Command(32'd70201404);
PIM_Command(32'd70401085);
PIM_Command(32'd87175998);
PIM_Command(32'd86980415);
PIM_Command(32'd87702336);
PIM_Command(32'd87111745);
PIM_Command(32'd87899714);
PIM_Command(32'd88097347);
PIM_Command(32'd88031556);
PIM_Command(32'd88031301);
PIM_Command(32'd88162886);
PIM_Command(32'd88359751);
PIM_Command(32'd71701832);
PIM_Command(32'd71435849);
PIM_Command(32'd71373898);
PIM_Command(32'd71636555);
PIM_Command(32'd71305292);
PIM_Command(32'd71241293);
PIM_Command(32'd71571534);
PIM_Command(32'd71767887);
PIM_Command(32'd71502160);
PIM_Command(32'd71699025);
PIM_Command(32'd71434322);
PIM_Command(32'd71370579);
PIM_Command(32'd71633748);
PIM_Command(32'd71303509);
PIM_Command(32'd71241558);
PIM_Command(32'd71566167);
PIM_Command(32'd71766104);
PIM_Command(32'd71500377);
PIM_Command(32'd89020250);
PIM_Command(32'd89412955);
PIM_Command(32'd89151580);
PIM_Command(32'd88689757);
PIM_Command(32'd88756830);
PIM_Command(32'd88624479);
PIM_Command(32'd88823392);
PIM_Command(32'd89807713);
PIM_Command(32'd88887138);
PIM_Command(32'd89217379);
PIM_Command(32'd89349732);
PIM_Command(32'd89808229);
PIM_Command(32'd88623718);
PIM_Command(32'd88821095);
PIM_Command(32'd88823912);
PIM_Command(32'd89150825);
PIM_Command(32'd89347946);
PIM_Command(32'd89414763);
PIM_Command(32'd89743212);
PIM_Command(32'd89939309);
PIM_Command(32'd90071150);
PIM_Command(32'd89940335);
PIM_Command(32'd90268272);
PIM_Command(32'd90136945);
PIM_Command(32'd90203250);
PIM_Command(32'd90400115);
PIM_Command(32'd90467444);
PIM_Command(32'd90534517);
PIM_Command(32'd90795638);
PIM_Command(32'd90664863);
PIM_Command(32'd91453086);
PIM_Command(32'd90928541);
PIM_Command(32'd90599324);
PIM_Command(32'd91255963);
PIM_Command(32'd91058586);
PIM_Command(32'd90730649);
PIM_Command(32'd90401432);
PIM_Command(32'd94872576);
PIM_Command(32'd296133633);
PIM_Command(32'd296199682);
PIM_Command(32'd94675715);
PIM_Command(32'd295936004);
PIM_Command(32'd94478341);
PIM_Command(32'd296091654);
PIM_Command(32'd83952903);
PIM_Command(32'd295699208);
PIM_Command(32'd84018185);
PIM_Command(32'd84018442);
PIM_Command(32'd84083979);
PIM_Command(32'd296026892);
PIM_Command(32'd94806285);
PIM_Command(32'd296027918);
PIM_Command(32'd84151567);
PIM_Command(32'd94570000);
PIM_Command(32'd296067601);
PIM_Command(32'd295870738);
PIM_Command(32'd296067859);
PIM_Command(32'd94834964);
PIM_Command(32'd83955989);
PIM_Command(32'd84742934);
PIM_Command(32'd84087319);
PIM_Command(32'd84481816);
PIM_Command(32'd84480537);
PIM_Command(32'd84612634);
PIM_Command(32'd67769627);
PIM_Command(32'd67110428);
PIM_Command(32'd85531421);
PIM_Command(32'd67572766);
PIM_Command(32'd85859103);
PIM_Command(32'd67835424);
PIM_Command(32'd67176481);
PIM_Command(32'd85598242);
PIM_Command(32'd68095523);
PIM_Command(32'd86188068);
PIM_Command(32'd67311653);
PIM_Command(32'd68163366);
PIM_Command(32'd86385959);
PIM_Command(32'd67242280);
PIM_Command(32'd86517033);
PIM_Command(32'd85793834);
PIM_Command(32'd85918763);
PIM_Command(32'd86122796);
PIM_Command(32'd86255917);
PIM_Command(32'd86648622);
PIM_Command(32'd86714671);
PIM_Command(32'd86779696);
PIM_Command(32'd86838321);
PIM_Command(32'd87044402);
PIM_Command(32'd70266419);
PIM_Command(32'd86979380);
PIM_Command(32'd86912821);
PIM_Command(32'd87110454);
PIM_Command(32'd70661431);
PIM_Command(32'd70529592);
PIM_Command(32'd70136121);
PIM_Command(32'd70596922);
PIM_Command(32'd87372603);
PIM_Command(32'd70201404);
PIM_Command(32'd70401085);
PIM_Command(32'd87175998);
PIM_Command(32'd86980415);
PIM_Command(32'd87702336);
PIM_Command(32'd87111745);
PIM_Command(32'd87899714);
PIM_Command(32'd88097347);
PIM_Command(32'd88031556);
PIM_Command(32'd88031301);
PIM_Command(32'd88162886);
PIM_Command(32'd88359751);
PIM_Command(32'd71701832);
PIM_Command(32'd71435849);
PIM_Command(32'd71373898);
PIM_Command(32'd71636555);
PIM_Command(32'd71305292);
PIM_Command(32'd71241293);
PIM_Command(32'd71571534);
PIM_Command(32'd71767887);
PIM_Command(32'd71502160);
PIM_Command(32'd71699025);
PIM_Command(32'd71434322);
PIM_Command(32'd71370579);
PIM_Command(32'd71633748);
PIM_Command(32'd71303509);
PIM_Command(32'd71241558);
PIM_Command(32'd71566167);
PIM_Command(32'd71766104);
PIM_Command(32'd71500377);
PIM_Command(32'd89020250);
PIM_Command(32'd89412955);
PIM_Command(32'd89151580);
PIM_Command(32'd88689757);
PIM_Command(32'd88756830);
PIM_Command(32'd88624479);
PIM_Command(32'd88823392);
PIM_Command(32'd89807713);
PIM_Command(32'd88887138);
PIM_Command(32'd89217379);
PIM_Command(32'd89349732);
PIM_Command(32'd89808229);
PIM_Command(32'd88623718);
PIM_Command(32'd88821095);
PIM_Command(32'd88823912);
PIM_Command(32'd89150825);
PIM_Command(32'd89347946);
PIM_Command(32'd89414763);
PIM_Command(32'd89743212);
PIM_Command(32'd89939309);
PIM_Command(32'd90071150);
PIM_Command(32'd89940335);
PIM_Command(32'd90268272);
PIM_Command(32'd90136945);
PIM_Command(32'd90203250);
PIM_Command(32'd90400115);
PIM_Command(32'd90467444);
PIM_Command(32'd90534517);
PIM_Command(32'd90795638);
PIM_Command(32'd90664871);
PIM_Command(32'd91453094);
PIM_Command(32'd90928549);
PIM_Command(32'd90599332);
PIM_Command(32'd91255971);
PIM_Command(32'd91058594);
PIM_Command(32'd90730657);
PIM_Command(32'd90401440);
PIM_Command(32'd95398912);
PIM_Command(32'd296659969);
PIM_Command(32'd296726018);
PIM_Command(32'd95202051);
PIM_Command(32'd296462340);
PIM_Command(32'd95004677);
PIM_Command(32'd296615942);
PIM_Command(32'd83952903);
PIM_Command(32'd296223496);
PIM_Command(32'd84018185);
PIM_Command(32'd84018442);
PIM_Command(32'd84083979);
PIM_Command(32'd296551180);
PIM_Command(32'd95332621);
PIM_Command(32'd296552206);
PIM_Command(32'd84151567);
PIM_Command(32'd95094288);
PIM_Command(32'd296593937);
PIM_Command(32'd296397074);
PIM_Command(32'd296594195);
PIM_Command(32'd95359252);
PIM_Command(32'd83955989);
PIM_Command(32'd84742934);
PIM_Command(32'd84087319);
PIM_Command(32'd84481816);
PIM_Command(32'd84480537);
PIM_Command(32'd84612634);
PIM_Command(32'd67769627);
PIM_Command(32'd67110428);
PIM_Command(32'd85531421);
PIM_Command(32'd67572766);
PIM_Command(32'd85859103);
PIM_Command(32'd67835424);
PIM_Command(32'd67176481);
PIM_Command(32'd85598242);
PIM_Command(32'd68095523);
PIM_Command(32'd86188068);
PIM_Command(32'd67311653);
PIM_Command(32'd68163366);
PIM_Command(32'd86385959);
PIM_Command(32'd67242280);
PIM_Command(32'd86517033);
PIM_Command(32'd85793834);
PIM_Command(32'd85918763);
PIM_Command(32'd86122796);
PIM_Command(32'd86255917);
PIM_Command(32'd86648622);
PIM_Command(32'd86714671);
PIM_Command(32'd86779696);
PIM_Command(32'd86838321);
PIM_Command(32'd87044402);
PIM_Command(32'd70266419);
PIM_Command(32'd86979380);
PIM_Command(32'd86912821);
PIM_Command(32'd87110454);
PIM_Command(32'd70661431);
PIM_Command(32'd70529592);
PIM_Command(32'd70136121);
PIM_Command(32'd70596922);
PIM_Command(32'd87372603);
PIM_Command(32'd70201404);
PIM_Command(32'd70401085);
PIM_Command(32'd87175998);
PIM_Command(32'd86980415);
PIM_Command(32'd87702336);
PIM_Command(32'd87111745);
PIM_Command(32'd87899714);
PIM_Command(32'd88097347);
PIM_Command(32'd88031556);
PIM_Command(32'd88031301);
PIM_Command(32'd88162886);
PIM_Command(32'd88359751);
PIM_Command(32'd71701832);
PIM_Command(32'd71435849);
PIM_Command(32'd71373898);
PIM_Command(32'd71636555);
PIM_Command(32'd71305292);
PIM_Command(32'd71241293);
PIM_Command(32'd71571534);
PIM_Command(32'd71767887);
PIM_Command(32'd71502160);
PIM_Command(32'd71699025);
PIM_Command(32'd71434322);
PIM_Command(32'd71370579);
PIM_Command(32'd71633748);
PIM_Command(32'd71303509);
PIM_Command(32'd71241558);
PIM_Command(32'd71566167);
PIM_Command(32'd71766104);
PIM_Command(32'd71500377);
PIM_Command(32'd89020250);
PIM_Command(32'd89412955);
PIM_Command(32'd89151580);
PIM_Command(32'd88689757);
PIM_Command(32'd88756830);
PIM_Command(32'd88624479);
PIM_Command(32'd88823392);
PIM_Command(32'd89807713);
PIM_Command(32'd88887138);
PIM_Command(32'd89217379);
PIM_Command(32'd89349732);
PIM_Command(32'd89808229);
PIM_Command(32'd88623718);
PIM_Command(32'd88821095);
PIM_Command(32'd88823912);
PIM_Command(32'd89150825);
PIM_Command(32'd89347946);
PIM_Command(32'd89414763);
PIM_Command(32'd89743212);
PIM_Command(32'd89939309);
PIM_Command(32'd90071150);
PIM_Command(32'd89940335);
PIM_Command(32'd90268272);
PIM_Command(32'd90136945);
PIM_Command(32'd90203250);
PIM_Command(32'd90400115);
PIM_Command(32'd90467444);
PIM_Command(32'd90534517);
PIM_Command(32'd90795638);
PIM_Command(32'd90664879);
PIM_Command(32'd91453102);
PIM_Command(32'd90928557);
PIM_Command(32'd90599340);
PIM_Command(32'd91255979);
PIM_Command(32'd91058602);
PIM_Command(32'd90730665);
PIM_Command(32'd90401448);
PIM_Command(32'd95925248);
PIM_Command(32'd297186305);
PIM_Command(32'd297252354);
PIM_Command(32'd95728387);
PIM_Command(32'd296988676);
PIM_Command(32'd95531013);
PIM_Command(32'd297140230);
PIM_Command(32'd83952903);
PIM_Command(32'd296747784);
PIM_Command(32'd84018185);
PIM_Command(32'd84018442);
PIM_Command(32'd84083979);
PIM_Command(32'd297075468);
PIM_Command(32'd95858957);
PIM_Command(32'd297076494);
PIM_Command(32'd84151567);
PIM_Command(32'd95618576);
PIM_Command(32'd297120273);
PIM_Command(32'd296923410);
PIM_Command(32'd297120531);
PIM_Command(32'd95883540);
PIM_Command(32'd83955989);
PIM_Command(32'd84742934);
PIM_Command(32'd84087319);
PIM_Command(32'd84481816);
PIM_Command(32'd84480537);
PIM_Command(32'd84612634);
PIM_Command(32'd67769627);
PIM_Command(32'd67110428);
PIM_Command(32'd85531421);
PIM_Command(32'd67572766);
PIM_Command(32'd85859103);
PIM_Command(32'd67835424);
PIM_Command(32'd67176481);
PIM_Command(32'd85598242);
PIM_Command(32'd68095523);
PIM_Command(32'd86188068);
PIM_Command(32'd67311653);
PIM_Command(32'd68163366);
PIM_Command(32'd86385959);
PIM_Command(32'd67242280);
PIM_Command(32'd86517033);
PIM_Command(32'd85793834);
PIM_Command(32'd85918763);
PIM_Command(32'd86122796);
PIM_Command(32'd86255917);
PIM_Command(32'd86648622);
PIM_Command(32'd86714671);
PIM_Command(32'd86779696);
PIM_Command(32'd86838321);
PIM_Command(32'd87044402);
PIM_Command(32'd70266419);
PIM_Command(32'd86979380);
PIM_Command(32'd86912821);
PIM_Command(32'd87110454);
PIM_Command(32'd70661431);
PIM_Command(32'd70529592);
PIM_Command(32'd70136121);
PIM_Command(32'd70596922);
PIM_Command(32'd87372603);
PIM_Command(32'd70201404);
PIM_Command(32'd70401085);
PIM_Command(32'd87175998);
PIM_Command(32'd86980415);
PIM_Command(32'd87702336);
PIM_Command(32'd87111745);
PIM_Command(32'd87899714);
PIM_Command(32'd88097347);
PIM_Command(32'd88031556);
PIM_Command(32'd88031301);
PIM_Command(32'd88162886);
PIM_Command(32'd88359751);
PIM_Command(32'd71701832);
PIM_Command(32'd71435849);
PIM_Command(32'd71373898);
PIM_Command(32'd71636555);
PIM_Command(32'd71305292);
PIM_Command(32'd71241293);
PIM_Command(32'd71571534);
PIM_Command(32'd71767887);
PIM_Command(32'd71502160);
PIM_Command(32'd71699025);
PIM_Command(32'd71434322);
PIM_Command(32'd71370579);
PIM_Command(32'd71633748);
PIM_Command(32'd71303509);
PIM_Command(32'd71241558);
PIM_Command(32'd71566167);
PIM_Command(32'd71766104);
PIM_Command(32'd71500377);
PIM_Command(32'd89020250);
PIM_Command(32'd89412955);
PIM_Command(32'd89151580);
PIM_Command(32'd88689757);
PIM_Command(32'd88756830);
PIM_Command(32'd88624479);
PIM_Command(32'd88823392);
PIM_Command(32'd89807713);
PIM_Command(32'd88887138);
PIM_Command(32'd89217379);
PIM_Command(32'd89349732);
PIM_Command(32'd89808229);
PIM_Command(32'd88623718);
PIM_Command(32'd88821095);
PIM_Command(32'd88823912);
PIM_Command(32'd89150825);
PIM_Command(32'd89347946);
PIM_Command(32'd89414763);
PIM_Command(32'd89743212);
PIM_Command(32'd89939309);
PIM_Command(32'd90071150);
PIM_Command(32'd89940335);
PIM_Command(32'd90268272);
PIM_Command(32'd90136945);
PIM_Command(32'd90203250);
PIM_Command(32'd90400115);
PIM_Command(32'd90467444);
PIM_Command(32'd90534517);
PIM_Command(32'd90795638);
PIM_Command(32'd90664887);
PIM_Command(32'd91453110);
PIM_Command(32'd90928565);
PIM_Command(32'd90599348);
PIM_Command(32'd91255987);
PIM_Command(32'd91058610);
PIM_Command(32'd90730673);
PIM_Command(32'd90401456);
PIM_Command(32'd96451584);
PIM_Command(32'd297712641);
PIM_Command(32'd297778690);
PIM_Command(32'd96254723);
PIM_Command(32'd297515012);
PIM_Command(32'd96057349);
PIM_Command(32'd297664518);
PIM_Command(32'd83952903);
PIM_Command(32'd297272072);
PIM_Command(32'd84018185);
PIM_Command(32'd84018442);
PIM_Command(32'd84083979);
PIM_Command(32'd297599756);
PIM_Command(32'd96385293);
PIM_Command(32'd297600782);
PIM_Command(32'd84151567);
PIM_Command(32'd96142864);
PIM_Command(32'd297646609);
PIM_Command(32'd297449746);
PIM_Command(32'd297646867);
PIM_Command(32'd96407828);
PIM_Command(32'd83955989);
PIM_Command(32'd84742934);
PIM_Command(32'd84087319);
PIM_Command(32'd84481816);
PIM_Command(32'd84480537);
PIM_Command(32'd84612634);
PIM_Command(32'd67769627);
PIM_Command(32'd67110428);
PIM_Command(32'd85531421);
PIM_Command(32'd67572766);
PIM_Command(32'd85859103);
PIM_Command(32'd67835424);
PIM_Command(32'd67176481);
PIM_Command(32'd85598242);
PIM_Command(32'd68095523);
PIM_Command(32'd86188068);
PIM_Command(32'd67311653);
PIM_Command(32'd68163366);
PIM_Command(32'd86385959);
PIM_Command(32'd67242280);
PIM_Command(32'd86517033);
PIM_Command(32'd85793834);
PIM_Command(32'd85918763);
PIM_Command(32'd86122796);
PIM_Command(32'd86255917);
PIM_Command(32'd86648622);
PIM_Command(32'd86714671);
PIM_Command(32'd86779696);
PIM_Command(32'd86838321);
PIM_Command(32'd87044402);
PIM_Command(32'd70266419);
PIM_Command(32'd86979380);
PIM_Command(32'd86912821);
PIM_Command(32'd87110454);
PIM_Command(32'd70661431);
PIM_Command(32'd70529592);
PIM_Command(32'd70136121);
PIM_Command(32'd70596922);
PIM_Command(32'd87372603);
PIM_Command(32'd70201404);
PIM_Command(32'd70401085);
PIM_Command(32'd87175998);
PIM_Command(32'd86980415);
PIM_Command(32'd87702336);
PIM_Command(32'd87111745);
PIM_Command(32'd87899714);
PIM_Command(32'd88097347);
PIM_Command(32'd88031556);
PIM_Command(32'd88031301);
PIM_Command(32'd88162886);
PIM_Command(32'd88359751);
PIM_Command(32'd71701832);
PIM_Command(32'd71435849);
PIM_Command(32'd71373898);
PIM_Command(32'd71636555);
PIM_Command(32'd71305292);
PIM_Command(32'd71241293);
PIM_Command(32'd71571534);
PIM_Command(32'd71767887);
PIM_Command(32'd71502160);
PIM_Command(32'd71699025);
PIM_Command(32'd71434322);
PIM_Command(32'd71370579);
PIM_Command(32'd71633748);
PIM_Command(32'd71303509);
PIM_Command(32'd71241558);
PIM_Command(32'd71566167);
PIM_Command(32'd71766104);
PIM_Command(32'd71500377);
PIM_Command(32'd89020250);
PIM_Command(32'd89412955);
PIM_Command(32'd89151580);
PIM_Command(32'd88689757);
PIM_Command(32'd88756830);
PIM_Command(32'd88624479);
PIM_Command(32'd88823392);
PIM_Command(32'd89807713);
PIM_Command(32'd88887138);
PIM_Command(32'd89217379);
PIM_Command(32'd89349732);
PIM_Command(32'd89808229);
PIM_Command(32'd88623718);
PIM_Command(32'd88821095);
PIM_Command(32'd88823912);
PIM_Command(32'd89150825);
PIM_Command(32'd89347946);
PIM_Command(32'd89414763);
PIM_Command(32'd89743212);
PIM_Command(32'd89939309);
PIM_Command(32'd90071150);
PIM_Command(32'd89940335);
PIM_Command(32'd90268272);
PIM_Command(32'd90136945);
PIM_Command(32'd90203250);
PIM_Command(32'd90400115);
PIM_Command(32'd90467444);
PIM_Command(32'd90534517);
PIM_Command(32'd90795638);
PIM_Command(32'd90664895);
PIM_Command(32'd91453118);
PIM_Command(32'd90928573);
PIM_Command(32'd90599356);
PIM_Command(32'd91255995);
PIM_Command(32'd91058618);
PIM_Command(32'd90730681);
PIM_Command(32'd90401464);
PIM_Command(32'd96977920);
PIM_Command(32'd298238977);
PIM_Command(32'd298305026);
PIM_Command(32'd96781059);
PIM_Command(32'd298041348);
PIM_Command(32'd96583685);
PIM_Command(32'd298188806);
PIM_Command(32'd83952903);
PIM_Command(32'd297796360);
PIM_Command(32'd84018185);
PIM_Command(32'd84018442);
PIM_Command(32'd84083979);
PIM_Command(32'd298124044);
PIM_Command(32'd96911629);
PIM_Command(32'd298125070);
PIM_Command(32'd84151567);
PIM_Command(32'd96667152);
PIM_Command(32'd298172945);
PIM_Command(32'd297976082);
PIM_Command(32'd298173203);
PIM_Command(32'd96932116);
PIM_Command(32'd83955989);
PIM_Command(32'd84742934);
PIM_Command(32'd84087319);
PIM_Command(32'd84481816);
PIM_Command(32'd84480537);
PIM_Command(32'd84612634);
PIM_Command(32'd67769627);
PIM_Command(32'd67110428);
PIM_Command(32'd85531421);
PIM_Command(32'd67572766);
PIM_Command(32'd85859103);
PIM_Command(32'd67835424);
PIM_Command(32'd67176481);
PIM_Command(32'd85598242);
PIM_Command(32'd68095523);
PIM_Command(32'd86188068);
PIM_Command(32'd67311653);
PIM_Command(32'd68163366);
PIM_Command(32'd86385959);
PIM_Command(32'd67242280);
PIM_Command(32'd86517033);
PIM_Command(32'd85793834);
PIM_Command(32'd85918763);
PIM_Command(32'd86122796);
PIM_Command(32'd86255917);
PIM_Command(32'd86648622);
PIM_Command(32'd86714671);
PIM_Command(32'd86779696);
PIM_Command(32'd86838321);
PIM_Command(32'd87044402);
PIM_Command(32'd70266419);
PIM_Command(32'd86979380);
PIM_Command(32'd86912821);
PIM_Command(32'd87110454);
PIM_Command(32'd70661431);
PIM_Command(32'd70529592);
PIM_Command(32'd70136121);
PIM_Command(32'd70596922);
PIM_Command(32'd87372603);
PIM_Command(32'd70201404);
PIM_Command(32'd70401085);
PIM_Command(32'd87175998);
PIM_Command(32'd86980415);
PIM_Command(32'd87702336);
PIM_Command(32'd87111745);
PIM_Command(32'd87899714);
PIM_Command(32'd88097347);
PIM_Command(32'd88031556);
PIM_Command(32'd88031301);
PIM_Command(32'd88162886);
PIM_Command(32'd88359751);
PIM_Command(32'd71701832);
PIM_Command(32'd71435849);
PIM_Command(32'd71373898);
PIM_Command(32'd71636555);
PIM_Command(32'd71305292);
PIM_Command(32'd71241293);
PIM_Command(32'd71571534);
PIM_Command(32'd71767887);
PIM_Command(32'd71502160);
PIM_Command(32'd71699025);
PIM_Command(32'd71434322);
PIM_Command(32'd71370579);
PIM_Command(32'd71633748);
PIM_Command(32'd71303509);
PIM_Command(32'd71241558);
PIM_Command(32'd71566167);
PIM_Command(32'd71766104);
PIM_Command(32'd71500377);
PIM_Command(32'd89020250);
PIM_Command(32'd89412955);
PIM_Command(32'd89151580);
PIM_Command(32'd88689757);
PIM_Command(32'd88756830);
PIM_Command(32'd88624479);
PIM_Command(32'd88823392);
PIM_Command(32'd89807713);
PIM_Command(32'd88887138);
PIM_Command(32'd89217379);
PIM_Command(32'd89349732);
PIM_Command(32'd89808229);
PIM_Command(32'd88623718);
PIM_Command(32'd88821095);
PIM_Command(32'd88823912);
PIM_Command(32'd89150825);
PIM_Command(32'd89347946);
PIM_Command(32'd89414763);
PIM_Command(32'd89743212);
PIM_Command(32'd89939309);
PIM_Command(32'd90071150);
PIM_Command(32'd89940335);
PIM_Command(32'd90268272);
PIM_Command(32'd90136945);
PIM_Command(32'd90203250);
PIM_Command(32'd90400115);
PIM_Command(32'd90467444);
PIM_Command(32'd90534517);
PIM_Command(32'd90795638);
PIM_Command(32'd90664903);
PIM_Command(32'd91453126);
PIM_Command(32'd90928581);
PIM_Command(32'd90599364);
PIM_Command(32'd91256003);
PIM_Command(32'd91058626);
PIM_Command(32'd90730689);
PIM_Command(32'd90401472);
PIM_Command(32'd97504256);
PIM_Command(32'd298765313);
PIM_Command(32'd298831362);
PIM_Command(32'd97307395);
PIM_Command(32'd298567684);
PIM_Command(32'd97110021);
PIM_Command(32'd298713094);
PIM_Command(32'd83952903);
PIM_Command(32'd298320648);
PIM_Command(32'd84018185);
PIM_Command(32'd84018442);
PIM_Command(32'd84083979);
PIM_Command(32'd298648332);
PIM_Command(32'd97437965);
PIM_Command(32'd298649358);
PIM_Command(32'd84151567);
PIM_Command(32'd97191440);
PIM_Command(32'd298699281);
PIM_Command(32'd298502418);
PIM_Command(32'd298699539);
PIM_Command(32'd97456404);
PIM_Command(32'd83955989);
PIM_Command(32'd84742934);
PIM_Command(32'd84087319);
PIM_Command(32'd84481816);
PIM_Command(32'd84480537);
PIM_Command(32'd84612634);
PIM_Command(32'd67769627);
PIM_Command(32'd67110428);
PIM_Command(32'd85531421);
PIM_Command(32'd67572766);
PIM_Command(32'd85859103);
PIM_Command(32'd67835424);
PIM_Command(32'd67176481);
PIM_Command(32'd85598242);
PIM_Command(32'd68095523);
PIM_Command(32'd86188068);
PIM_Command(32'd67311653);
PIM_Command(32'd68163366);
PIM_Command(32'd86385959);
PIM_Command(32'd67242280);
PIM_Command(32'd86517033);
PIM_Command(32'd85793834);
PIM_Command(32'd85918763);
PIM_Command(32'd86122796);
PIM_Command(32'd86255917);
PIM_Command(32'd86648622);
PIM_Command(32'd86714671);
PIM_Command(32'd86779696);
PIM_Command(32'd86838321);
PIM_Command(32'd87044402);
PIM_Command(32'd70266419);
PIM_Command(32'd86979380);
PIM_Command(32'd86912821);
PIM_Command(32'd87110454);
PIM_Command(32'd70661431);
PIM_Command(32'd70529592);
PIM_Command(32'd70136121);
PIM_Command(32'd70596922);
PIM_Command(32'd87372603);
PIM_Command(32'd70201404);
PIM_Command(32'd70401085);
PIM_Command(32'd87175998);
PIM_Command(32'd86980415);
PIM_Command(32'd87702336);
PIM_Command(32'd87111745);
PIM_Command(32'd87899714);
PIM_Command(32'd88097347);
PIM_Command(32'd88031556);
PIM_Command(32'd88031301);
PIM_Command(32'd88162886);
PIM_Command(32'd88359751);
PIM_Command(32'd71701832);
PIM_Command(32'd71435849);
PIM_Command(32'd71373898);
PIM_Command(32'd71636555);
PIM_Command(32'd71305292);
PIM_Command(32'd71241293);
PIM_Command(32'd71571534);
PIM_Command(32'd71767887);
PIM_Command(32'd71502160);
PIM_Command(32'd71699025);
PIM_Command(32'd71434322);
PIM_Command(32'd71370579);
PIM_Command(32'd71633748);
PIM_Command(32'd71303509);
PIM_Command(32'd71241558);
PIM_Command(32'd71566167);
PIM_Command(32'd71766104);
PIM_Command(32'd71500377);
PIM_Command(32'd89020250);
PIM_Command(32'd89412955);
PIM_Command(32'd89151580);
PIM_Command(32'd88689757);
PIM_Command(32'd88756830);
PIM_Command(32'd88624479);
PIM_Command(32'd88823392);
PIM_Command(32'd89807713);
PIM_Command(32'd88887138);
PIM_Command(32'd89217379);
PIM_Command(32'd89349732);
PIM_Command(32'd89808229);
PIM_Command(32'd88623718);
PIM_Command(32'd88821095);
PIM_Command(32'd88823912);
PIM_Command(32'd89150825);
PIM_Command(32'd89347946);
PIM_Command(32'd89414763);
PIM_Command(32'd89743212);
PIM_Command(32'd89939309);
PIM_Command(32'd90071150);
PIM_Command(32'd89940335);
PIM_Command(32'd90268272);
PIM_Command(32'd90136945);
PIM_Command(32'd90203250);
PIM_Command(32'd90400115);
PIM_Command(32'd90467444);
PIM_Command(32'd90534517);
PIM_Command(32'd90795638);
PIM_Command(32'd90664911);
PIM_Command(32'd91453134);
PIM_Command(32'd90928589);
PIM_Command(32'd90599372);
PIM_Command(32'd91256011);
PIM_Command(32'd91058634);
PIM_Command(32'd90730697);
PIM_Command(32'd90401480);
PIM_Command(32'd98030592);
PIM_Command(32'd299291649);
PIM_Command(32'd299357698);
PIM_Command(32'd97833731);
PIM_Command(32'd299094020);
PIM_Command(32'd97636357);
PIM_Command(32'd299237382);
PIM_Command(32'd83952903);
PIM_Command(32'd298844936);
PIM_Command(32'd84018185);
PIM_Command(32'd84018442);
PIM_Command(32'd84083979);
PIM_Command(32'd299172620);
PIM_Command(32'd97964301);
PIM_Command(32'd299173646);
PIM_Command(32'd84151567);
PIM_Command(32'd97715728);
PIM_Command(32'd299225617);
PIM_Command(32'd299028754);
PIM_Command(32'd299225875);
PIM_Command(32'd97980692);
PIM_Command(32'd83955989);
PIM_Command(32'd84742934);
PIM_Command(32'd84087319);
PIM_Command(32'd84481816);
PIM_Command(32'd84480537);
PIM_Command(32'd84612634);
PIM_Command(32'd67769627);
PIM_Command(32'd67110428);
PIM_Command(32'd85531421);
PIM_Command(32'd67572766);
PIM_Command(32'd85859103);
PIM_Command(32'd67835424);
PIM_Command(32'd67176481);
PIM_Command(32'd85598242);
PIM_Command(32'd68095523);
PIM_Command(32'd86188068);
PIM_Command(32'd67311653);
PIM_Command(32'd68163366);
PIM_Command(32'd86385959);
PIM_Command(32'd67242280);
PIM_Command(32'd86517033);
PIM_Command(32'd85793834);
PIM_Command(32'd85918763);
PIM_Command(32'd86122796);
PIM_Command(32'd86255917);
PIM_Command(32'd86648622);
PIM_Command(32'd86714671);
PIM_Command(32'd86779696);
PIM_Command(32'd86838321);
PIM_Command(32'd87044402);
PIM_Command(32'd70266419);
PIM_Command(32'd86979380);
PIM_Command(32'd86912821);
PIM_Command(32'd87110454);
PIM_Command(32'd70661431);
PIM_Command(32'd70529592);
PIM_Command(32'd70136121);
PIM_Command(32'd70596922);
PIM_Command(32'd87372603);
PIM_Command(32'd70201404);
PIM_Command(32'd70401085);
PIM_Command(32'd87175998);
PIM_Command(32'd86980415);
PIM_Command(32'd87702336);
PIM_Command(32'd87111745);
PIM_Command(32'd87899714);
PIM_Command(32'd88097347);
PIM_Command(32'd88031556);
PIM_Command(32'd88031301);
PIM_Command(32'd88162886);
PIM_Command(32'd88359751);
PIM_Command(32'd71701832);
PIM_Command(32'd71435849);
PIM_Command(32'd71373898);
PIM_Command(32'd71636555);
PIM_Command(32'd71305292);
PIM_Command(32'd71241293);
PIM_Command(32'd71571534);
PIM_Command(32'd71767887);
PIM_Command(32'd71502160);
PIM_Command(32'd71699025);
PIM_Command(32'd71434322);
PIM_Command(32'd71370579);
PIM_Command(32'd71633748);
PIM_Command(32'd71303509);
PIM_Command(32'd71241558);
PIM_Command(32'd71566167);
PIM_Command(32'd71766104);
PIM_Command(32'd71500377);
PIM_Command(32'd89020250);
PIM_Command(32'd89412955);
PIM_Command(32'd89151580);
PIM_Command(32'd88689757);
PIM_Command(32'd88756830);
PIM_Command(32'd88624479);
PIM_Command(32'd88823392);
PIM_Command(32'd89807713);
PIM_Command(32'd88887138);
PIM_Command(32'd89217379);
PIM_Command(32'd89349732);
PIM_Command(32'd89808229);
PIM_Command(32'd88623718);
PIM_Command(32'd88821095);
PIM_Command(32'd88823912);
PIM_Command(32'd89150825);
PIM_Command(32'd89347946);
PIM_Command(32'd89414763);
PIM_Command(32'd89743212);
PIM_Command(32'd89939309);
PIM_Command(32'd90071150);
PIM_Command(32'd89940335);
PIM_Command(32'd90268272);
PIM_Command(32'd90136945);
PIM_Command(32'd90203250);
PIM_Command(32'd90400115);
PIM_Command(32'd90467444);
PIM_Command(32'd90534517);
PIM_Command(32'd90795638);
PIM_Command(32'd90664919);
PIM_Command(32'd91453142);
PIM_Command(32'd90928597);
PIM_Command(32'd90599380);
PIM_Command(32'd91256019);
PIM_Command(32'd91058642);
PIM_Command(32'd90730705);
PIM_Command(32'd90401488);
PIM_Command(32'd98556928);
PIM_Command(32'd299817985);
PIM_Command(32'd299884034);
PIM_Command(32'd98360067);
PIM_Command(32'd299620356);
PIM_Command(32'd98162693);
PIM_Command(32'd299761670);
PIM_Command(32'd83952903);
PIM_Command(32'd299369224);
PIM_Command(32'd84018185);
PIM_Command(32'd84018442);
PIM_Command(32'd84083979);
PIM_Command(32'd299696908);
PIM_Command(32'd98490637);
PIM_Command(32'd299697934);
PIM_Command(32'd84151567);
PIM_Command(32'd98240016);
PIM_Command(32'd299751953);
PIM_Command(32'd299555090);
PIM_Command(32'd299752211);
PIM_Command(32'd98504980);
PIM_Command(32'd83955989);
PIM_Command(32'd84742934);
PIM_Command(32'd84087319);
PIM_Command(32'd84481816);
PIM_Command(32'd84480537);
PIM_Command(32'd84612634);
PIM_Command(32'd67769627);
PIM_Command(32'd67110428);
PIM_Command(32'd85531421);
PIM_Command(32'd67572766);
PIM_Command(32'd85859103);
PIM_Command(32'd67835424);
PIM_Command(32'd67176481);
PIM_Command(32'd85598242);
PIM_Command(32'd68095523);
PIM_Command(32'd86188068);
PIM_Command(32'd67311653);
PIM_Command(32'd68163366);
PIM_Command(32'd86385959);
PIM_Command(32'd67242280);
PIM_Command(32'd86517033);
PIM_Command(32'd85793834);
PIM_Command(32'd85918763);
PIM_Command(32'd86122796);
PIM_Command(32'd86255917);
PIM_Command(32'd86648622);
PIM_Command(32'd86714671);
PIM_Command(32'd86779696);
PIM_Command(32'd86838321);
PIM_Command(32'd87044402);
PIM_Command(32'd70266419);
PIM_Command(32'd86979380);
PIM_Command(32'd86912821);
PIM_Command(32'd87110454);
PIM_Command(32'd70661431);
PIM_Command(32'd70529592);
PIM_Command(32'd70136121);
PIM_Command(32'd70596922);
PIM_Command(32'd87372603);
PIM_Command(32'd70201404);
PIM_Command(32'd70401085);
PIM_Command(32'd87175998);
PIM_Command(32'd86980415);
PIM_Command(32'd87702336);
PIM_Command(32'd87111745);
PIM_Command(32'd87899714);
PIM_Command(32'd88097347);
PIM_Command(32'd88031556);
PIM_Command(32'd88031301);
PIM_Command(32'd88162886);
PIM_Command(32'd88359751);
PIM_Command(32'd71701832);
PIM_Command(32'd71435849);
PIM_Command(32'd71373898);
PIM_Command(32'd71636555);
PIM_Command(32'd71305292);
PIM_Command(32'd71241293);
PIM_Command(32'd71571534);
PIM_Command(32'd71767887);
PIM_Command(32'd71502160);
PIM_Command(32'd71699025);
PIM_Command(32'd71434322);
PIM_Command(32'd71370579);
PIM_Command(32'd71633748);
PIM_Command(32'd71303509);
PIM_Command(32'd71241558);
PIM_Command(32'd71566167);
PIM_Command(32'd71766104);
PIM_Command(32'd71500377);
PIM_Command(32'd89020250);
PIM_Command(32'd89412955);
PIM_Command(32'd89151580);
PIM_Command(32'd88689757);
PIM_Command(32'd88756830);
PIM_Command(32'd88624479);
PIM_Command(32'd88823392);
PIM_Command(32'd89807713);
PIM_Command(32'd88887138);
PIM_Command(32'd89217379);
PIM_Command(32'd89349732);
PIM_Command(32'd89808229);
PIM_Command(32'd88623718);
PIM_Command(32'd88821095);
PIM_Command(32'd88823912);
PIM_Command(32'd89150825);
PIM_Command(32'd89347946);
PIM_Command(32'd89414763);
PIM_Command(32'd89743212);
PIM_Command(32'd89939309);
PIM_Command(32'd90071150);
PIM_Command(32'd89940335);
PIM_Command(32'd90268272);
PIM_Command(32'd90136945);
PIM_Command(32'd90203250);
PIM_Command(32'd90400115);
PIM_Command(32'd90467444);
PIM_Command(32'd90534517);
PIM_Command(32'd90795638);
PIM_Command(32'd90664927);
PIM_Command(32'd91453150);
PIM_Command(32'd90928605);
PIM_Command(32'd90599388);
PIM_Command(32'd91256027);
PIM_Command(32'd91058650);
PIM_Command(32'd90730713);
PIM_Command(32'd90401496);
PIM_Command(32'd99083264);
PIM_Command(32'd300344321);
PIM_Command(32'd300410370);
PIM_Command(32'd98886403);
PIM_Command(32'd300146692);
PIM_Command(32'd98689029);
PIM_Command(32'd300285958);
PIM_Command(32'd83952903);
PIM_Command(32'd299893512);
PIM_Command(32'd84018185);
PIM_Command(32'd84018442);
PIM_Command(32'd84083979);
PIM_Command(32'd300221196);
PIM_Command(32'd99016973);
PIM_Command(32'd300222222);
PIM_Command(32'd84151567);
PIM_Command(32'd98764304);
PIM_Command(32'd300278289);
PIM_Command(32'd300081426);
PIM_Command(32'd300278547);
PIM_Command(32'd99029268);
PIM_Command(32'd83955989);
PIM_Command(32'd84742934);
PIM_Command(32'd84087319);
PIM_Command(32'd84481816);
PIM_Command(32'd84480537);
PIM_Command(32'd84612634);
PIM_Command(32'd67769627);
PIM_Command(32'd67110428);
PIM_Command(32'd85531421);
PIM_Command(32'd67572766);
PIM_Command(32'd85859103);
PIM_Command(32'd67835424);
PIM_Command(32'd67176481);
PIM_Command(32'd85598242);
PIM_Command(32'd68095523);
PIM_Command(32'd86188068);
PIM_Command(32'd67311653);
PIM_Command(32'd68163366);
PIM_Command(32'd86385959);
PIM_Command(32'd67242280);
PIM_Command(32'd86517033);
PIM_Command(32'd85793834);
PIM_Command(32'd85918763);
PIM_Command(32'd86122796);
PIM_Command(32'd86255917);
PIM_Command(32'd86648622);
PIM_Command(32'd86714671);
PIM_Command(32'd86779696);
PIM_Command(32'd86838321);
PIM_Command(32'd87044402);
PIM_Command(32'd70266419);
PIM_Command(32'd86979380);
PIM_Command(32'd86912821);
PIM_Command(32'd87110454);
PIM_Command(32'd70661431);
PIM_Command(32'd70529592);
PIM_Command(32'd70136121);
PIM_Command(32'd70596922);
PIM_Command(32'd87372603);
PIM_Command(32'd70201404);
PIM_Command(32'd70401085);
PIM_Command(32'd87175998);
PIM_Command(32'd86980415);
PIM_Command(32'd87702336);
PIM_Command(32'd87111745);
PIM_Command(32'd87899714);
PIM_Command(32'd88097347);
PIM_Command(32'd88031556);
PIM_Command(32'd88031301);
PIM_Command(32'd88162886);
PIM_Command(32'd88359751);
PIM_Command(32'd71701832);
PIM_Command(32'd71435849);
PIM_Command(32'd71373898);
PIM_Command(32'd71636555);
PIM_Command(32'd71305292);
PIM_Command(32'd71241293);
PIM_Command(32'd71571534);
PIM_Command(32'd71767887);
PIM_Command(32'd71502160);
PIM_Command(32'd71699025);
PIM_Command(32'd71434322);
PIM_Command(32'd71370579);
PIM_Command(32'd71633748);
PIM_Command(32'd71303509);
PIM_Command(32'd71241558);
PIM_Command(32'd71566167);
PIM_Command(32'd71766104);
PIM_Command(32'd71500377);
PIM_Command(32'd89020250);
PIM_Command(32'd89412955);
PIM_Command(32'd89151580);
PIM_Command(32'd88689757);
PIM_Command(32'd88756830);
PIM_Command(32'd88624479);
PIM_Command(32'd88823392);
PIM_Command(32'd89807713);
PIM_Command(32'd88887138);
PIM_Command(32'd89217379);
PIM_Command(32'd89349732);
PIM_Command(32'd89808229);
PIM_Command(32'd88623718);
PIM_Command(32'd88821095);
PIM_Command(32'd88823912);
PIM_Command(32'd89150825);
PIM_Command(32'd89347946);
PIM_Command(32'd89414763);
PIM_Command(32'd89743212);
PIM_Command(32'd89939309);
PIM_Command(32'd90071150);
PIM_Command(32'd89940335);
PIM_Command(32'd90268272);
PIM_Command(32'd90136945);
PIM_Command(32'd90203250);
PIM_Command(32'd90400115);
PIM_Command(32'd90467444);
PIM_Command(32'd90534517);
PIM_Command(32'd90795638);
PIM_Command(32'd90664935);
PIM_Command(32'd91453158);
PIM_Command(32'd90928613);
PIM_Command(32'd90599396);
PIM_Command(32'd91256035);
PIM_Command(32'd91058658);
PIM_Command(32'd90730721);
PIM_Command(32'd90401504);
PIM_Command(32'd99609600);
PIM_Command(32'd300870657);
PIM_Command(32'd300936706);
PIM_Command(32'd99412739);
PIM_Command(32'd300673028);
PIM_Command(32'd99215365);
PIM_Command(32'd300810246);
PIM_Command(32'd83952903);
PIM_Command(32'd300417800);
PIM_Command(32'd84018185);
PIM_Command(32'd84018442);
PIM_Command(32'd84083979);
PIM_Command(32'd300745484);
PIM_Command(32'd99543309);
PIM_Command(32'd300746510);
PIM_Command(32'd84151567);
PIM_Command(32'd99288592);
PIM_Command(32'd300804625);
PIM_Command(32'd300607762);
PIM_Command(32'd300804883);
PIM_Command(32'd99553556);
PIM_Command(32'd83955989);
PIM_Command(32'd84742934);
PIM_Command(32'd84087319);
PIM_Command(32'd84481816);
PIM_Command(32'd84480537);
PIM_Command(32'd84612634);
PIM_Command(32'd67769627);
PIM_Command(32'd67110428);
PIM_Command(32'd85531421);
PIM_Command(32'd67572766);
PIM_Command(32'd85859103);
PIM_Command(32'd67835424);
PIM_Command(32'd67176481);
PIM_Command(32'd85598242);
PIM_Command(32'd68095523);
PIM_Command(32'd86188068);
PIM_Command(32'd67311653);
PIM_Command(32'd68163366);
PIM_Command(32'd86385959);
PIM_Command(32'd67242280);
PIM_Command(32'd86517033);
PIM_Command(32'd85793834);
PIM_Command(32'd85918763);
PIM_Command(32'd86122796);
PIM_Command(32'd86255917);
PIM_Command(32'd86648622);
PIM_Command(32'd86714671);
PIM_Command(32'd86779696);
PIM_Command(32'd86838321);
PIM_Command(32'd87044402);
PIM_Command(32'd70266419);
PIM_Command(32'd86979380);
PIM_Command(32'd86912821);
PIM_Command(32'd87110454);
PIM_Command(32'd70661431);
PIM_Command(32'd70529592);
PIM_Command(32'd70136121);
PIM_Command(32'd70596922);
PIM_Command(32'd87372603);
PIM_Command(32'd70201404);
PIM_Command(32'd70401085);
PIM_Command(32'd87175998);
PIM_Command(32'd86980415);
PIM_Command(32'd87702336);
PIM_Command(32'd87111745);
PIM_Command(32'd87899714);
PIM_Command(32'd88097347);
PIM_Command(32'd88031556);
PIM_Command(32'd88031301);
PIM_Command(32'd88162886);
PIM_Command(32'd88359751);
PIM_Command(32'd71701832);
PIM_Command(32'd71435849);
PIM_Command(32'd71373898);
PIM_Command(32'd71636555);
PIM_Command(32'd71305292);
PIM_Command(32'd71241293);
PIM_Command(32'd71571534);
PIM_Command(32'd71767887);
PIM_Command(32'd71502160);
PIM_Command(32'd71699025);
PIM_Command(32'd71434322);
PIM_Command(32'd71370579);
PIM_Command(32'd71633748);
PIM_Command(32'd71303509);
PIM_Command(32'd71241558);
PIM_Command(32'd71566167);
PIM_Command(32'd71766104);
PIM_Command(32'd71500377);
PIM_Command(32'd89020250);
PIM_Command(32'd89412955);
PIM_Command(32'd89151580);
PIM_Command(32'd88689757);
PIM_Command(32'd88756830);
PIM_Command(32'd88624479);
PIM_Command(32'd88823392);
PIM_Command(32'd89807713);
PIM_Command(32'd88887138);
PIM_Command(32'd89217379);
PIM_Command(32'd89349732);
PIM_Command(32'd89808229);
PIM_Command(32'd88623718);
PIM_Command(32'd88821095);
PIM_Command(32'd88823912);
PIM_Command(32'd89150825);
PIM_Command(32'd89347946);
PIM_Command(32'd89414763);
PIM_Command(32'd89743212);
PIM_Command(32'd89939309);
PIM_Command(32'd90071150);
PIM_Command(32'd89940335);
PIM_Command(32'd90268272);
PIM_Command(32'd90136945);
PIM_Command(32'd90203250);
PIM_Command(32'd90400115);
PIM_Command(32'd90467444);
PIM_Command(32'd90534517);
PIM_Command(32'd90795638);
PIM_Command(32'd90664943);
PIM_Command(32'd91453166);
PIM_Command(32'd90928621);
PIM_Command(32'd90599404);
PIM_Command(32'd91256043);
PIM_Command(32'd91058666);
PIM_Command(32'd90730729);
PIM_Command(32'd90401512);
PIM_Command(32'd100135936);
PIM_Command(32'd301396993);
PIM_Command(32'd301463042);
PIM_Command(32'd99939075);
PIM_Command(32'd301199364);
PIM_Command(32'd99741701);
PIM_Command(32'd301334534);
PIM_Command(32'd83952903);
PIM_Command(32'd300942088);
PIM_Command(32'd84018185);
PIM_Command(32'd84018442);
PIM_Command(32'd84083979);
PIM_Command(32'd301269772);
PIM_Command(32'd100069645);
PIM_Command(32'd301270798);
PIM_Command(32'd84151567);
PIM_Command(32'd99812880);
PIM_Command(32'd301330961);
PIM_Command(32'd301134098);
PIM_Command(32'd301331219);
PIM_Command(32'd100077844);
PIM_Command(32'd83955989);
PIM_Command(32'd84742934);
PIM_Command(32'd84087319);
PIM_Command(32'd84481816);
PIM_Command(32'd84480537);
PIM_Command(32'd84612634);
PIM_Command(32'd67769627);
PIM_Command(32'd67110428);
PIM_Command(32'd85531421);
PIM_Command(32'd67572766);
PIM_Command(32'd85859103);
PIM_Command(32'd67835424);
PIM_Command(32'd67176481);
PIM_Command(32'd85598242);
PIM_Command(32'd68095523);
PIM_Command(32'd86188068);
PIM_Command(32'd67311653);
PIM_Command(32'd68163366);
PIM_Command(32'd86385959);
PIM_Command(32'd67242280);
PIM_Command(32'd86517033);
PIM_Command(32'd85793834);
PIM_Command(32'd85918763);
PIM_Command(32'd86122796);
PIM_Command(32'd86255917);
PIM_Command(32'd86648622);
PIM_Command(32'd86714671);
PIM_Command(32'd86779696);
PIM_Command(32'd86838321);
PIM_Command(32'd87044402);
PIM_Command(32'd70266419);
PIM_Command(32'd86979380);
PIM_Command(32'd86912821);
PIM_Command(32'd87110454);
PIM_Command(32'd70661431);
PIM_Command(32'd70529592);
PIM_Command(32'd70136121);
PIM_Command(32'd70596922);
PIM_Command(32'd87372603);
PIM_Command(32'd70201404);
PIM_Command(32'd70401085);
PIM_Command(32'd87175998);
PIM_Command(32'd86980415);
PIM_Command(32'd87702336);
PIM_Command(32'd87111745);
PIM_Command(32'd87899714);
PIM_Command(32'd88097347);
PIM_Command(32'd88031556);
PIM_Command(32'd88031301);
PIM_Command(32'd88162886);
PIM_Command(32'd88359751);
PIM_Command(32'd71701832);
PIM_Command(32'd71435849);
PIM_Command(32'd71373898);
PIM_Command(32'd71636555);
PIM_Command(32'd71305292);
PIM_Command(32'd71241293);
PIM_Command(32'd71571534);
PIM_Command(32'd71767887);
PIM_Command(32'd71502160);
PIM_Command(32'd71699025);
PIM_Command(32'd71434322);
PIM_Command(32'd71370579);
PIM_Command(32'd71633748);
PIM_Command(32'd71303509);
PIM_Command(32'd71241558);
PIM_Command(32'd71566167);
PIM_Command(32'd71766104);
PIM_Command(32'd71500377);
PIM_Command(32'd89020250);
PIM_Command(32'd89412955);
PIM_Command(32'd89151580);
PIM_Command(32'd88689757);
PIM_Command(32'd88756830);
PIM_Command(32'd88624479);
PIM_Command(32'd88823392);
PIM_Command(32'd89807713);
PIM_Command(32'd88887138);
PIM_Command(32'd89217379);
PIM_Command(32'd89349732);
PIM_Command(32'd89808229);
PIM_Command(32'd88623718);
PIM_Command(32'd88821095);
PIM_Command(32'd88823912);
PIM_Command(32'd89150825);
PIM_Command(32'd89347946);
PIM_Command(32'd89414763);
PIM_Command(32'd89743212);
PIM_Command(32'd89939309);
PIM_Command(32'd90071150);
PIM_Command(32'd89940335);
PIM_Command(32'd90268272);
PIM_Command(32'd90136945);
PIM_Command(32'd90203250);
PIM_Command(32'd90400115);
PIM_Command(32'd90467444);
PIM_Command(32'd90534517);
PIM_Command(32'd90795638);
PIM_Command(32'd90664951);
PIM_Command(32'd91453174);
PIM_Command(32'd90928629);
PIM_Command(32'd90599412);
PIM_Command(32'd91256051);
PIM_Command(32'd91058674);
PIM_Command(32'd90730737);
PIM_Command(32'd90401520);
PIM_Command(32'd100662272);
PIM_Command(32'd301923329);
PIM_Command(32'd301989378);
PIM_Command(32'd100465411);
PIM_Command(32'd301725700);
PIM_Command(32'd100268037);
PIM_Command(32'd301858822);
PIM_Command(32'd83952903);
PIM_Command(32'd301466376);
PIM_Command(32'd84018185);
PIM_Command(32'd84018442);
PIM_Command(32'd84083979);
PIM_Command(32'd301794060);
PIM_Command(32'd100595981);
PIM_Command(32'd301795086);
PIM_Command(32'd84151567);
PIM_Command(32'd100337168);
PIM_Command(32'd301857297);
PIM_Command(32'd301660434);
PIM_Command(32'd301857555);
PIM_Command(32'd100602132);
PIM_Command(32'd83955989);
PIM_Command(32'd84742934);
PIM_Command(32'd84087319);
PIM_Command(32'd84481816);
PIM_Command(32'd84480537);
PIM_Command(32'd84612634);
PIM_Command(32'd67769627);
PIM_Command(32'd67110428);
PIM_Command(32'd85531421);
PIM_Command(32'd67572766);
PIM_Command(32'd85859103);
PIM_Command(32'd67835424);
PIM_Command(32'd67176481);
PIM_Command(32'd85598242);
PIM_Command(32'd68095523);
PIM_Command(32'd86188068);
PIM_Command(32'd67311653);
PIM_Command(32'd68163366);
PIM_Command(32'd86385959);
PIM_Command(32'd67242280);
PIM_Command(32'd86517033);
PIM_Command(32'd85793834);
PIM_Command(32'd85918763);
PIM_Command(32'd86122796);
PIM_Command(32'd86255917);
PIM_Command(32'd86648622);
PIM_Command(32'd86714671);
PIM_Command(32'd86779696);
PIM_Command(32'd86838321);
PIM_Command(32'd87044402);
PIM_Command(32'd70266419);
PIM_Command(32'd86979380);
PIM_Command(32'd86912821);
PIM_Command(32'd87110454);
PIM_Command(32'd70661431);
PIM_Command(32'd70529592);
PIM_Command(32'd70136121);
PIM_Command(32'd70596922);
PIM_Command(32'd87372603);
PIM_Command(32'd70201404);
PIM_Command(32'd70401085);
PIM_Command(32'd87175998);
PIM_Command(32'd86980415);
PIM_Command(32'd87702336);
PIM_Command(32'd87111745);
PIM_Command(32'd87899714);
PIM_Command(32'd88097347);
PIM_Command(32'd88031556);
PIM_Command(32'd88031301);
PIM_Command(32'd88162886);
PIM_Command(32'd88359751);
PIM_Command(32'd71701832);
PIM_Command(32'd71435849);
PIM_Command(32'd71373898);
PIM_Command(32'd71636555);
PIM_Command(32'd71305292);
PIM_Command(32'd71241293);
PIM_Command(32'd71571534);
PIM_Command(32'd71767887);
PIM_Command(32'd71502160);
PIM_Command(32'd71699025);
PIM_Command(32'd71434322);
PIM_Command(32'd71370579);
PIM_Command(32'd71633748);
PIM_Command(32'd71303509);
PIM_Command(32'd71241558);
PIM_Command(32'd71566167);
PIM_Command(32'd71766104);
PIM_Command(32'd71500377);
PIM_Command(32'd89020250);
PIM_Command(32'd89412955);
PIM_Command(32'd89151580);
PIM_Command(32'd88689757);
PIM_Command(32'd88756830);
PIM_Command(32'd88624479);
PIM_Command(32'd88823392);
PIM_Command(32'd89807713);
PIM_Command(32'd88887138);
PIM_Command(32'd89217379);
PIM_Command(32'd89349732);
PIM_Command(32'd89808229);
PIM_Command(32'd88623718);
PIM_Command(32'd88821095);
PIM_Command(32'd88823912);
PIM_Command(32'd89150825);
PIM_Command(32'd89347946);
PIM_Command(32'd89414763);
PIM_Command(32'd89743212);
PIM_Command(32'd89939309);
PIM_Command(32'd90071150);
PIM_Command(32'd89940335);
PIM_Command(32'd90268272);
PIM_Command(32'd90136945);
PIM_Command(32'd90203250);
PIM_Command(32'd90400115);
PIM_Command(32'd90467444);
PIM_Command(32'd90534517);
PIM_Command(32'd90795638);
PIM_Command(32'd90664959);
PIM_Command(32'd91453182);
PIM_Command(32'd90928637);
PIM_Command(32'd90599420);
PIM_Command(32'd91256059);
PIM_Command(32'd91058682);
PIM_Command(32'd90730745);
PIM_Command(32'd90401528);



endtask


endmodule