task test_simon();
    $display("SIMON Program");
endtask