task test_ecb_aes();
    $display("ECB AES Program");
endtask